��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�
�����@Xk���Fq���$Z�u�չ���J 	��Ǐ�J;a��^��?�o{̛������^���P�C����L�9jc��?3�8*���	̆����=H���Wݝ�QE���o��d)J�%����e���vid��:�x�y��d|W̱p�)^�MJ"y^.F��)�zg�����^yje�ӟ�:��:� @+�K�O�n�D JA���l(�Z2L�x�_)8Y�(��U�@iG��� �����-ix���L�DB6c^F~,$������FD��;�m�������!�������)J�:�w��8�����ȅ�|��������)
����ȪD���xkE�[,�D�n�)�t#�Ym���&����&
�u$����,~�j��C���j6��nI�ZEwd:�D�iT7��[����� ��/��ÔP�������m�={���l���F�y�����yI���s��_�R��mɜﻄ�_U���N�M��wr�1��
�7��!�U~_�4�Q��}j��vҦJ���4_z0���4꾻rM|`vW5����D�r�D�GX7xh{@+[�Yx�6͜�=��5?�،��qj�y�+�]���_>ĝ����'�&Խ򔱈��2i��P�V��&
!�>�r"5M$p#J��g,>�T��)ŀ6m��a~���m6V)�$܀2t@N�\"d�{�/';� ���T���b*j�����D�I;|��'�4���@ߨfz�+	8Y(�B��g�Mq�g�:��-D�RF厯�o�c.���)iO���n	V�Z�ay�xf�k$,��>Z[��/��������ar�6'�fG�<��S����G�³P����?b
�rB� ��t��u��L@�*�j�	Q��p/Ǡ�������l�8�����u'V�!���'0�>w9U�16J�H��P���ODA���n��6���<�G�����=i2��[���u�!��<�;����|(��"�R\7OW�Ѧ�y�v���" y����L ��8,J��X�4#I��{��)zD��;��+F\׵�sqE9`vl8^�Q?	����D,�Q��m<�oNxT����j�+g�������V�q��k1�ؗ�&�GwUs`�h^L{�����Lه��
�|�ߜm�(D�~$��wЬ���^�d]�����rW�7�d�b-M*#��}�>o�����Ղ~��*N���� ��������d�F��)�:ꈇ����"�,��f�0�p���u&cs�����ʯ�v���#b��%��'֪4�U���l Uc�q������Hh5�wX۰�)ݴ2��%�3c�("C�
e�nT9��$)$^�����V��J��WQ�~PC%!3r�ps�4e�p��V$'�|B�d>/k�=�<ڌ>j!A8o*��j;�Z�AF���͕�����[BU��gA����%@��K���w�v�>SӠ]���y)X��Q�檴7��|Jg����X���� 3��&��=���;-þ��f&�O78/��ȉ�L�[%=PDa��8��ǳ�ʿ�z%y:��R$Un~H����	3z�j�7�߾:I����f�'�0Vv�_EW�(�}�ۄ���ں'�]�
�f�Ǽ�._V7e5�G��=צr�UsE;��+����[s���z�*I��:�۪\��e������ھU��I�,?��ŗk�Z �!����r��:���
���(X�s%h��2�LbD��[Ǐ�f�HQ^" �����O�&����p)�A���](�^GKy��,�S\0,��y���fr��B``}�5�����f�=rT&�E\ݓ��'���n�b��א��|�U��QG�G�oU����ځ9�e.���h�n��H����=|����	����7���^�r!�o"�|�7�@�i8�E���~�EK��kҸ��ǘ3M�'q�,����PK�f�wC�X�)�y֊��iA�a�f��^S���f�iϧ�+��q� �M<ji1dZA����@�37���ո7��1����}��6�w�#���v�UKIzkf��!]\c���.�f <� �ű�픋/4�?�C$�n+��$0v��o��M��N@��Ƶ��f�+m�%o���$���M�ў�g6D��=�hSu^u+,�b���R�(�:�nڹ�y�FX6�Y�qL�����ܐkU �8�Ve�������ų@�?��Y��Ԡ�-5=6T�y����+Ve��"*���P���}�=/�g��m�/Zr�eU�v0���l���!����B*�
7����
X��.Ó�ޚ"x~�=���	GB��o�
���\�~�(s���<wo�&����|ި�u���2�l��}���s.������y�MS�qp�%�LY	�� B8 ޴��`Fj�q�M:���Z��:�_�V�-M��i�	��K�o
�C���c))���m�\w~�q��s�r�e������LlnS�{Y���[V�b�|{T�d���ճ�^�@z��;��V���!�O�{쇆�(e��.\����^���9ԘV�����҆س��c�O9����wi���y媀,	��t�/�_������G|��\w�� B]�D��u��9��4
�OY��� (N�>����N*!ޙܟ�Y�s�a��`�{�	[=�Z�0x!�%�hw�}i4"25_�u�n��/(p'�+ݳ���܊�Y�=��f�?�WJ)��x�SEey~ģD"�`�H���p���y���4&�����եad=���j����p0��a������UѮZ�0��i3��b�i��>�H��R�*��۴B��H�P��Sf�U0�O�:\�V�-�U��"���w���=@�v����sf��1+=��ס�U��	�!���{cv���W��'l߀j�k��ӿg�&&
	|ȡA kt��I�(%���=[��ZUl�w��3�Ƽ~�(���*'�s>�-Ń5r;`�I�ݦ&�]�v�I�~�1��o.`�Z%!�j{^ׇ��W��T�v2�E�CMn��	5p*�J�Q� �G�\�]��N���jˑ��`K��$Sm�Z�^FY�����ߊ�o5Y f�7W����Nj���,?o=��MG�O��b���K;���cW,��b"ǺI���}������ds�[�~�����a�*b�yQl����kd��a��;�1%�V&x���JQ.J�/����������IˤQȾ�Oy���J8�q$��Ezh�O5#�9�;�.��c^Mam�c�쀜����:C��0'���>�3l�����)�Y�ۭIu�����$�6���#�
�V:BJ!pt�L���=s�b6xA�����!��glbP�p ��>�7ս�ق�
�XU�c�]�)��D����ND����RR0��C{�*���x�*�:a���R$�����!@@H��3��z�	]%�Fo��
_e����;6m4�x�E4N�D�NFn�7~Z#ȭ��ڒ�������U!ˠ��웙,�b�p����� ���En̾J��t�>5�qm6�p�I�e���}W������'s��Wi����ú���s׶��w�G_��Z_a��@���O���ɯ�7߃��U��gy\q>_IE�g;���Ϳ�:f)�Y���[b�n[�ȫ C�SPWVȤ��]e���Z�S��>PͿ�6�>d���<��~�J�Zcg��B�:���{����؜z��4�5��ផ11���O[l��(O��_��5���L����I<����]�k[똎� ��O�`nN������<�a���E�ym<�뀒eh��*(/��a̭1s����X��	�CkY�:�^���A`mVT�7��/VtMo���1�L~Q��=���v0ԬC���[w*/v*��Jm]&��g�h��u./^��}v�~)����p�FG��A�H����דڙ��/���Af����-u�\��(|��+0���\}��)LT�އ�&N�	S����?!sI�B�B����s�.I�l� �Φ�G+��`���c����$n%)�+BK�1Oh�I	��
Iz#:
�5/Q��;�Q�?�ٟ�nV�{$�Mc:C<)�%�*�=�އpU*e�U�^�n��Ӆ��S��38�;Nț~Gf1Sfҽ��<k��[Nu >��~�oR�3"�Sv.ϋ���%�����hC���5�ʫuy>Hhj�%RݘK�&��X��'4�k�FA��ߨ��V�nsr�3'�^BR'2~�V!����e �s@1��,�@�tR��0MZ��� �5��=t�=|�&��_��H��U�??�[�K���㉆1�a`�&
T{{���)\Jۘ�f��f"�r�Ѩ� ��ϫ8%C���1ݕF�o�X�戔>P.|(����Ŧ�JF�6������cr�H����d`V\\��[��)��YJ!� �*![co��a�����7ֲ��B�eF�����.�kɎn����{Q8�/���%H������~E��ˀ�X�Ժ�N�O��W�C��l�h:N�[����O��/=k����WV�_%��{�qP'��Qo�/�jF����g{3m��J������7b�D�%��ĦN���l��&�^�j�+_��ky�99c�>�&Xb������k�&$�+��`�sK��3�đ�3�����(�$ݙ�D�q5$� h�i�Io:�c��*��=:�K�z�rMn��^�����&.�F�0�d�OI9{M�����M. �O�}휥����QG�1=>�!p��)�[�(����[����0�E��|ȇF���ʷf�
2�ֵ>c�`�2d5���h�� �~�3�\;H}���r��������C�'��N�~���o�}�� <+گ�ǈ��Q]�٦t�f1�v��Pg�2�lh��Z�(�5]]���5��sN���4_!{�I=��F㓱�pن���s���j��+�͍e�v�e�$�=��P=��q�K h��R�o��d���&��o(q{�\�U��A��o%�TV���JLxc�#ʣJWɵu�(�WR劄ň�7�)��Vw�QX����_�Y%7��;������'E��@۲ H��j'm�~nup�m<���������_�<d�f��	nb�?F~��60��B��Ԉ^	�>�
9�T�����N��+�g��͜���!ޭ��5���t�ٵ��涻��f�
B��h\���Ė ���_��z	�W��?�t���V�:����z���C�߀��p~��yg��w�V��aa�7	e �����@��s�g���
t}����z��-��ώ�i�:��O4����FPB�!$H\��hater�g�KX?��gH#|�Ps�]K��Ձ�ڟ�	$�&����p��evn��_���-�4N�Z,$y��r�9摇�]wA��y���z�c�Vz )@�+�7M�qk"@�}�%�,�-+��7o#F\��̽w�5�w����r,�����Ɨ~{�������U9Bdy+�I���J|��.���L!�=�8��F��/u_<�<"q�:!�!�_��}�G?�)��;(��W��-�v�mE� ��}�Di���+�97�1T����3гo���9R�t��${�p��d?��ڑ"#Zy�'����'��!��tbM����R1,pkB�f
Z�Z9�s�Ϧ��z�*��;�ʤ�b5+Cz��u>���Rlw
�0�Tfd��!�'��9�Is��\g7_\�����o��JRs�U�/P����?h[���^�G=-XZ�*R��}�q��	�����ϴ�{(����'����`+:��[{����aS􁾨H�	�n����o�E�:��t�6&�É�.�l��IF1�m�]���[A�w9rZ�-�b���'=�I_w��dK']ܷ3
�|6�����U��j4]�Mp��ӌ�ZT���:t'���ѱ+EȢ�~8%.%�nA{��F�b[[���4V�[��h�b��I"�s�Cc�2��U�Gx�HF�G��
�����3��{`�Վ�v������=����IE�T?02h��l�h�P�;\��� �݂��O���ɗFt�Cr鍪��a8T�Dq��E��������j'&�����hf���=2r;w �������TdjR ���MH��c��7ȜlF�R���l��Q�M����0��_��p�H\��;v��-è��k�!��#�+55�-. �QF[h�Iݡ�-�=瘎��3$���=
�뜈��G��q�@�.�=M���GI¨�eT[h��O!��'���r�}���q�d�ok��9 ᯀ$�:�9|�e���_�.:�Pq@ӵH�|gQ̫�E��g�'k0:x#d���"0�=�-�
�,G��c�ٖ4A��Ǻd��?8^�_T�W����¶J��-2ߟ��P�Í ���� b�$k7\��wC�zV)`�y��e�ܥ�@�5��:;NB�E��;�qn) m/�mˮj8ǱcB�4�����gb ]�S�0"5�8�a���/u�QT%��z�f鑔�y���h��
J=���?�Ѱ�KrI�[�2�����g�8��)���z+]2�/�~�	��6�ƅ%�4{)[���ˇ~OQRr�[���_m�xvD�4�t��x���������X"y&�Mt8�[y��L{���5S� [��`�l8�=%r��P���_�Ϥ��Շ�0���
K6�3�*�F��7����e�}�~�Z������Ҕ��bz��
ha�µ�URO��|B�dC�z+�>k0��)��z6�A"�� ƽ�k���P)�0-���e�!���������g����K�4x��d/*���b�Z��Sp+-Y��>��B�ӌ��z]џS%a�j��n\��x��!&�k+��%�az�`��)��DRT%ܲE�K蚸���H9#��zP���;uY��"9���87"W�7A5��|�r��ktї�����Լb��0�$��i? L�1!����.�DO
(����SE#��%}v��W-9M�0�� � �e���z���y��7	�c���^ިW��6	ݗ���-,�a@5��w��w)d����1Ϛ�b�J�\I�T�?S@�0��U�.�*�K6�ׅ��b	TZ�̰&o�Lu����D�A��g�]?"�
��ʘ�\Е�]X�=�?��B��=@�z�Դ�>Ci�0`� *,�G���i����Nb��&�~	�M�%#��-�&@���w#g��)��]��0(p@�>W��Z�M���'{�+I��#���O1�;����6��D6��=N�.�>����JR��L�� ��Ρ@���?���J1	7�_|�挭�PãK���T�*9�DU0������wI��'a�W�F-����O�l<�Z��Ú�j��è���XY�,�A'O�Y�`���Ά����TV1� �3�]jԬ�UC�k,3*�D"�Z��j\\C\���}�;�Yvķ�mn�"���i�V�.�<�z"�.1��0:7n����FZ���}� �5Nn����*�KŤm=B�ʃָ�T0��	�[BWHQ�A��
̆���	hӘ���i�Ѻ��t;F*��s5(j3�10FI��!�g95��O�o��%y߱�b��#A@|��귾���x{�h�>�DJ�gt��*�K�gv�V]_�GW!�ˈ'�Wj�]{ ����{�5�J͎�]õ��sAI��+3�_t��"�L��43K���& <�ׯas�����
ؾ4]2?�y���0y~�T���W�8�0c2f/=:t��p�\��'�\�(���&�w!v��-ޏ�~�%꙼#��������3��J/�U-��o���{�+#�bگ��Eߧ/m�H@�1pU��ׂ�p+�9#��+�0�G��%w�¥]ňP9�u'zw����
�r���"��B��"��Q];�g���r��`�C�h�	�J"�=����/��/�+�����'QbI�]�F�d��Ç��b
.�=��sS�E�ތ �dV����������LΗ�ˡ=m���E���(��G|��*��9I^I|�7���X./PӞ���E� ����CMۍ�{Ib��X�2��$���װH�U��Y�ڌ�����˃\s5����O� �c������=�`��-K
�:I��OK�Ex�_2�9 ��by4}���n�n&+� u��F�z�H�5.��])_D���^RP=��	����sfTC����a)z���	[�-���w2����{�1$0�a��|&�:���Q�F�"=�����o�:��Q�ث:cš�rLu�~�g	�-���8"��g��L1���<Ԛ���ϝ�X�ʯ{ٷ��­�b"�-ʖ�j?jp�3�p���0Ѵ�A��w@�⑨���o�����[CK�p�F����g��r9Uν��ʿ$	�x2�`��(��oQo���h�zk�C��V��������xi�u�^2��C({Ok�U��P�'��!ʁ�YO,d��j�%��5=�2�X/vm�*�,Ӹ%]�l+%O��"�p��w��o:�)@��/I�	p�WT^Z8���1�W)�,'(�[P	��1͡���G�B%cR����3f	�/f�ޝ���2	#5�!J���q�4�ev��yו.���#�3n��4�������A�"t&��|��?��EB����.�|X#xl
���%���+�΅2�F$1�4s���׍�\��Иv%o�P��_��4����ƪY3�Fb����徉?��-�	�a(~m!T���|(�f]��sW�V�J����R�����IН�׫�y�Y��7�x@�}�%p�_"?����
D�*#^I��0�H!����S���=�΅�F��Tw_�˝eY+���ZǍ���J�Պ^yOx���?�e*��(�wR�ώ/IG;��כ�Htp�*K����i�J/'D�d��2U�v:�k�i�v�]e�+F,�LI�Ug{���*'@�]�<�C����H��[�׶:�vCR6�K��;b��[��b!V���F+r>�5�Ǟ�PC�G�z�������QM����e���6��K�3iBI������^Y����O>:�Zp�ݼ��I��
��s�0�[r��@��ib�̒@˗HA��WG��v@���P�9��H��ƅ�+�,Gr@��~)²�
�؇
��3�\�5���i���Z��������p��+��:��b�X?:��ì�Ѓ^�l�(���EhP�#�0)]�ou+���ҥ�Ȝn���%gk�ϼ!�p�xn��i���)�ړ$9�E)���ot �q-�ps��`O��g��\�м����웓F~�$d$�6�W�@�����(��f��O�O���\�9]�)F��}KҖ��oQjY�R̃j�������-�j:4I �����"�^芘i��N�i~f��q�Z���+
Tr�f�@�u��-�V��h���D��T�`�Iv9��c�B��M�M�G���9�#kG�P�ϡ��k���8H_�$�c��0vM�2Μ�}wPb�ή�[�R;z��l��e�z�����@O{���#+��f��ik6�`5�f�Qq�1���O6�j�쐲@�;8����:��/�r*!��rB�(��X�c�)�w�\;Yz��lb@��7�a%-��O-��0��\⦂s־r�G�H�S�V� 0�|�����`]�$@P]�PL�a�x��_�3�(��?m�I����l��"�U��Q"�lJt"���WE;�������� �Ͽ��MVPP���;���ͯ:Jp�>H3k����V��y���N�mMMX�z�&1Z[��⯰���������z%ݓ��ebXl`w���f�_�(���h��#KHk�Ε;L���'~�I
���� F�3��dY��I��<^�=���"��-5�xx�p��=ʮu4}����T'R[����EO��uK��5m8���D)�Q��6��*YN��ӱ�·�4�S�����7I2�H�e.e�B���>^�
/�Z/�ˎ�\�ܡ�t��w��Ky@��k��*�ᮭ���pW�	�!���rF(�,p�o�� }o�u��WWd�f��p�]����б�4��`t�����^U���}r��SN�����a5]!`%��A~�%?�F�Ǭ'����~��^�X�e�[v�+p�j��0%NL��̎�ߎ��H+T==),X��/�i�Va��;�UF�)h��6�\��8�|���2�jXk��7��H���\�-�bh��Сz��m�{��_0H�x�z(�ީn�j�1��l��(�&3�V��D�QE������V�F�3.�4G��ԛ�@�h�è,@|��)~(��cS�+@�&Vg9�v	4�*�-]�b{[x %T����Щ5��_�p�;�u���'��c7�<;�k����M���H0�r�8��Wt p�E�Xji���&�"BW;�����*�a1oA�W�3 ��aGܮ����&�33kw��E'Zg4��sQ���P�pPu���\Yǃ���ox���� �_����UE�T���U�̍��i�:�����#���:W<��x�B�1m�Nn�^Պye��7�J���p���$��=~�t2�ɹ�����?!c��Y&��U��&�f.�G��;hr>(H��!����� ]LZR�x�Bω�t�Ơ>�U:$Mt� ��i����q�g�&!ke�:uD[�����y	 |�Ww�\�_	c����oo��H8�rwE��B�Ɉ�_���?�(�X#oC�z������g��1JOn�����Hm���kpZs(fLs+_%��#x�����`��ifx6���M�3ˈ#�;��[�#������Xx��6e�����aL&W-��,l��X����z�Ej�����ˌDIm��<� 53��Ԋ�er��*L��h>��U��	�ޭ8�-W;��O~�W���9e����d�d���	z[c9�b�c�!}(5���K�8`L��WE�b����X��$���즪����ۗw�Y��y^��~RDl�p�STМ�^�W��dm�6���%��}^�tU_�0c4��z/N�Z�}L?NE�Ln��F��'\��7�7t����*�����2ɚ�������@$�t<eVS�R�L,�-5�B��[��#�h�J���ҏ�%3&��
g�!��3c1Q^j����`{̧����H�y��h�����6��$��SpK�K�/��^gj�%	�F@Tm�<7�~��If4'TDJ|��	�Ntţ>�U���a�̷����;�K�,�A�j�����/nMW�بÚ�f�w��I^>ݰ���{t��P��;�g .?Æ ^L)��?z*Ņ��������q���	���ֹ��Р������qp����#�X�Q�IM$�����2ǝ�SCC-�Qq�TQA�t}ڪ
#��Z�Ma�/�?����r0s��p���"q�
��XS�b��F��� �h�����KJ�=��KglD*�����{7�hv˖�ր�:��guo�r�� ��v�ܬ�� �x�o��8a2��%�0��,�@D�5=�<��tչX����>9>NJ���},���2��J�C��D�}n`2�%-�X��,�@7%N�iwO��L�'\�����QR�2�_*X�m�S�ꃲ�U�uv~��-?�tB��p�w�M$U�k�}MV� : "������T�i��KS�J;�a@g��N�R������ς�%#���׼�"<C�r��ثEj����Ê�������8$-S�=h9{��9o$8TY�S �̝��ɮ��Ggf�����(8�#4),�I�Zo�0N�ń���Ea&8����S�;��3����["���j^��[Ek�Bi2� �bK��H'w@C_Y;,���<v���'@���/�a�r��m�̓�EӲ�
��b��	8R`F.	zO���?b�W.7qz�W�W<Eԁ�ҧ9h��g�)���@q1>�Q��g���$�P9���C�60(���X�=J��Uq�hD��3�
�ᱰq�C�2~�1�����ϥҼ&����#�s�<0�F)���#���K�^6�]���s���}�9y�����Y��]�&G�w�(��]��M쌰"-�������X� �Q~�D���OTH������&����p��n���>6Ty��aX���	C�1�T8��X�"�r�%�>^K�7Jb܃4y��[c��{����	�̟�q�?P�HL���;�)�������r��\��w��3���p������/��M�,�ׅ�����2l+�2��$	Z�ҫA� �+��I[�Q֗�F�G4=I0F���:�c�ַ���0�W�Jݒ�������ˠ_뤢9A��Ƞ�[n�T~2C�r���71����Q}�����ۈ�����q�`��1x�p��i�C��3����s��,�F�L�L��o��l���>�lH��ws��# �K3!y�>\�����}�¢��tb�[)6<KL��^�}?8�2yk��-6lRj�ńF���H5����J	y`�`ݭ7 ��nՒj�g��#�b���������a*H�F\�B֓�Q�'ö5��N�~��lQ=��{Q��Z���&U�u��T��g�EҒ��&�ʖ�C�y�(4GG��uL1ʦcq�m6=�`�G���8w�C�ݪ����Ԝm�&:�;�qT#�=e��	��+}����l
�k*E,x�o[Qt��\�������-����������>+�b�L���8L1��z�}>VW�7��,�@��/�=�F���
4 �R����#��~Q�5�ɚ�cw	��J����"�=
�b� B����:b��c���9Ս��,A
�٨1݀O�@�Q�b��Q���!@�������L
���Ըt���Ŝ(ъ���[�T�܏������#yV+���?#�v�CF�{����v���_(2o-����1�U�;���r��=�udMf��@^l�x��A�9ڦb)~b�BԶ@m$ t��	�HM��^z��e��@�-�M�}c6��������)�Lý�6�A��5��2l���Rod'��7��?F�bv"���'ƥ9*��{���N���.����o"��8|%���T���%N��L���l�ʑ{�z��m�P�9Oq�7k}0e���Cd�4�����w���Ja�8�M���ͻI2P��3�G5�8�-�OU��ݎ�]fH�-�"����&�I1>����w����KO�� t��o�������f�5�r��>�22�����*�1_X��n���K0�Lsu������z�_�l*_�45�� ��`�Y^�PZ��ǝR�K�Si�����b�:}�]TK�w�Zt�d~Q��`��F�Nx\������{"�NVy3BЉ$KS�ή/�J؏�����<���o!+�ymE(��ެ�RP����x��9�\�U���Q�����/5���Glz�T1%���}r;�� B��e�����*�"`�_Q�*p9��Y*��{�kOA�"��`'w�A�B7����&Sh�6��{�B�5��j���%"���:�o]܇�?�|v��6ω@X8��r����x��^9p��b���	��W��M�貾
��I�>����<�	�)_��Y .x�^/5A���0I^����&���V�>r�klw>�d�=NG�К.��	�D6��H��C�����m�d��Y��L�D�`��� :v�ӵ�E�*����Kt�
�b��9�f����]M�qb	X�G��h���Rи�;KRA�<V ��H��5�6��ԫ�0���v���N�?�%�y�9�i�n�Z5�,�G��_��-�Z��fkQ��a��۲n��UmYǷ�ض��/¢�m����#�s�f�?|W���@�4����k�9 9�D�1��)�I
���\\~&��ڡf�]���=��?LF	�3���貨���s�k9�'
� ��0�w�ڭ��d�'��,�	���8�&`�{�|�8%�Î:�I*z3��)�G��;c�W�K��љ�=AfS��I�!�elh����r�J�Ʀ��7���w�pJ�k�y�(`\M~�����ܩT?7W���n����}|���\���55�Y�YCPxI۽'�:�b�T|/^�v��M�C|��5tQ���8��SOz������Q�f�"M7�a��	�q�i*�\�ȽT[P{R,-�U�k-����vu��B��f5������{u,ׅ��*Y���O́�����+�ْ
`b#L`^�?a�3�����d�2�#��߲�*���ÍXE�����d8�1obǐ��s��ő��h�5d�x��|�1��T?��&�� ĝ�=崓?����^��ڢ[�ը���X'X(�e�_�x�rKbȮ\��k�����,���0!�
q��:�~Hn���Y����@W���dT�M���;�m Cim�/4���@ls����Bɠ���ڟo�?U�Sa��(? 9�)O�����a�m�j��B��LЎ�aQ�	��ݖY��fG� mȫo��1p�c2��ߏa�`�z����PD�+�&��$�n]�Μ�i=x�
C,xڈ��M!����͗��S�a���fO�[(b0@]�Y��F�E����B�3�,�  D���訒B����5_g^s�g̎[��)b���.���:���8��KrȽ��}n�V�1�����f�҂���L#_�k�LJ������k&i�,�l봟)*)�r��8�_�B��}8*�m��
�#�����s"�]���j���⚖��ׅ��Gkm��s�c	Od��˙�wW�s�qo-�l�����|?V����;���I���5��o������Y��\��u�*��Ci'��$v)������'����I|ZT�e�DDA�8ꇃ^q8;���N��X\0�U��=&á���Ǿ�_u����4fl��"x������;���!��	��xb[��B&5�R����G����)��������!�ðG��˝���L�yX
c U����5M�X7"-������!$���
��.�f��w����T�Dz$��Hx|B1�6"4�� K#��%�_���'!#7ۗśUG���'2:F�����j�����(�����X�s�⠈[�;����I�e�"�| ��)L�Il�F7�j�����fR��+�b�n�z��@l�$h7�Xٛ'�	Um
5�f�h���ꃙ��V�+�~���?�f�h�#c�ģ��~�Z��"�~B�0�T8�6�˗��DM�r�8���Ջ����׸��;UPȜR���iTcC�6V9�}�bt@���Εv��F}X�G�{O��ZaAu�79o��ZME�h��r*7�0�����!`pМ��8g��Ƨ���ȥy�8��pfȜۿ������ω���\��8t��t���ɑ����S!c�I92,�hH_��2��f�3��0�ZT$��h�}{V������o��3G��[l�
�ݑ�C45�#��[�G�>*�ڿԱ���*d���g�����n�ys-�JE���r��)��l�pߍn���+N�p�yw��e_)�S��z�z��1S֖�Æ�����
aib&vz��;�EtI�\B�M+>��,܁�Nd�~V�^hR77}��z�A��1�f:�I�)�P6��.��Ъ�*�ߝ��#+��!d�J�(�Fm�@�E�H�i�	����m�8M�*���l��|m�>.�޼�f�'5�q��UC�k�	2��������X�@�ج�����;*��������<n�g6g7��i��_�����=��uca@��멏�j�>��z1/qO[���	����dg�E�3n�K?s*[�]�G����z����g�q<�?/\���!��x5P� 1V?�}G���%���@���Ύo�c&�=�_�����|y�v4$]��qK�Ej޷��ﳧ��.�>���!��!V�Ji�53�/�h.�
>��a�sC���Z�_ �Y�����Xy&

�ˀ�+f��ϭ�	���H���Fr�v�1P ��[y����[`q [y��%L(Ʈ�ߖ"�x_���F��������u��z��c���nf"���/���e�Z�ؿ��)�ѡ˹1쩃�T��z]�&6�l�������[��+��8�܍���
lZ����eP��Q�0dXN.�7?�)���uXR��7��3��FAܳ��j�#%�C�	�.�j��eʷ�춁�o�E���?�ֲ�w�0s��Ψ$ջ����o�k���>�X�d�������H���P�H�������[Ċ"n:� ��E��6>��a�c��j$�@V���f��.�f��*B��i�U��~�
��_'!.��H�/��@���S]��A͋)}� :_���o�+�=�j("��- ]/�A���|�=h~��k��4ᘓf��&�8��h�������H0-�4��|�4;sRe�:[ �p������en��k�K�&�fwV(�\��ʆk��8j��a7�[��̓����ٟ<na�o�M�C ���L��]�j+���kp�xr3.�^K�=����Ci���g��9$�>�w@3�1�����pe� �R�����3�J%"a8'�mz��� �h4�}��#����<>���xf>Q7�(�_���S1�3!oL��r��F����WfS�9RJG�h
ֻs\d�As�PaY���&1�>,�h��a�;P���y;G�R���y��%=E�����!D}�oP���F��¨�>�O5�p�8Y�[ZK�	�:,m�q�56}mi{�1��ć�m�mؐ{�|i�N{������ @�"�{w�Sg��Bߪ -������r%I{0�i` �Z5*s!ɒM ]���o�1�/`c��H_vev���oΆ�k�ޮ�:!�i(�k�)��CL{�?��0���[����<�9R�|O��I�M����>�`�u�V�ޘn�LGoB���\��!���I݆�N�a�p�vO�Ә�cޭF	*��p;6��XI�W�O��P�U��|��
�Ax8Ӈ�Lyv��C1D��P�!��������d��g�03�lSq���O������Z'�1�.�"kVMd#NߘwI�P�|���S%l)�ku�-��	�imԋm�����lb�ʣ�-�cX��a�5�'_ ��OC0� Gݸ����1%��~W �S���l�Mz���3�������l��s��_;��͟L�ܐO�1;� ��"k��[�V� &�D?�ٝx��'	�R�H��#L���uq�G;:�,ᒯl�מ�Em=&��Q�ڏ���ґY
�f
��
�&��ä�?݇�
P�R�DUh�	��Ű��ʵ�F���h�42W���wtFE�9m�rV�`���r�6�d�{�"-��(ޡ)G�7Dxc��#��DHF�4�B��T�������(��W���zr�%�\ߦ�2]���Yg��W�v������x�n?SjՀ!�v^��$W��<g*���B���,lqY�v��q�и>�q3�����b5H7��Am�ɻ 	=����%_�.�6{ȼ�o�WO0YM�ORT�NN)�'��C���ܔ�;�z���Bʹ,g|s��%�p�T��"��3'������\�z)������!�G��1��ZF��������4L�U?�ac�7͜�9��8�Z!��莅x̝��Ђ�xY�}_�b!i��K���q[�mZcG���S�y�<��7`�
���<�r>��{_^�?��j�������~��t�Y��������|��][_��hΞjT�p��k��{��#N\��ӳm�t�eK�?=|���oL�����m��%;8�aAV���K����qæ�"h�� J?ȬZq)u�u*���f�F*��i�W�-��Q;��g@)�n/�ӄ�d�i|m��B�\��U����,''�(�{2�@=�+���7aoQ��;��۱�kP�	�I U��R��?����$�c�;��7��_��߶���>�+��?9)q����!'
Q}������?��__
:������C^��:hd�N.�Z��s-[���^ױ ߐև�5���-�c�bK}�!�u����`�q �s������q�Inf��u5
�#�}Q7�o��$�4Ղ����M)%�V��?L�
���W+m�Ys��
��e=���?��h8��D9�QZ�,��H�S� �̙8d���Ϡ�q��5�B"9�od�ĝ�_Ox��|��6�a�؞(w��qyd��3A�%�W�#�z]P��70 ��E���o�V�b��݌yS����Ѣg�����!��F'$&�w�f?%�V8��/�=r���ф��>H3�XG^ ��/�8ČN*��l�ѩP@�W���t��%�a�F��q�D��8gg�_[> D1N-��)aB�����j��vGN�ʖ=�v�j߈p����L|�b���\ܫ��8O�-
����I�RH�� s
�`�'Lx�i��V��h�p�䨅���?����
�ɷԞ�C7Þ�S��KRf��([���+;��Ҕ�P�vs&fe<��D�m�ѹ������k�y��q?�$���Z�4b�z�{����@
�Ǌ�� &`�� 1���˸/!|]q<o&���h�ؗ�(4!������f�Y�\�&B�����蹷$/�qz<�+�T�,h���-���TA�aD5������/IPz�W���VS,�ж:���soi����R�|L�FW�c���c@d��S�̴���P	m%�t�~P��������BuI�dB:ŉc��u�e����O	l`�i��<�ۤ���n�}����Q��T��P��
�f�ubP𡧔lMYϬ >��F:��Y���yF�_:����g]�� ����i���r����\����R�;4��M����-��{���V<�[Y���������$}Ȝ�ox8�0��q)f���:5'�`�7R��<���(�ʵln"��-;�F�x�i^�	��:�l�BS˿y;O��W�6R��z������¥d�G��U���!�a�� ������[�8�"�u	pR��=3��IHS�c�Ƙ�cUXђ��PEv�ח�������tty��U�6
?2I��	�ڐ�kQu!X��Dۓ��,�_ޱ*3[Y���ߕ��E�!�6�� m*7���M�6�e�D�QC#�؄����L��,+.n/ʻL��(P�#�d؉J��TOz1>����e ����&�휬�s�o�x-)�p!��I�Ք���+6��JG�:V5PIr�j����[�,����m��4�G�����V�C�
}
RZc�*�[�uy���o5	���K�e�ۛ�S�劜4lf�G����>���q�z���1212��C�*���|~6q�&P��q�9 ��r�;��=��)?꠮eO�a#ն�օ؝|=k���u��.�i����4�\�M�L5���q��aiヾ��5��+ݜ'/�����pk�s�Q(3!@�8U��d?!<o! �:�_냮�
v���_~����֐ۏ� 	��u��y��C<H��`&����d�����A�	4���M����C� ���#�
Z�Q��JI�������#tF�߯`�
�Ql�{�<�<�b����u���}�3%0��$ϱ�7��#<���w^d�8��"�f�|f�8l��f��Є���{��M�&�vs��"Є���Q3���Iw;�&fûo�5���ABN���IP���O�EV��Iuɟ!"��̥�ݯ�/��6��È�j�p6D}�����e&6?�y��Fc���f��rn��N�%$��R8L��k��w��G�j���Pb�U����#ЫF�lƏs���������;�w�6�چM���4\zс� /a��k{#Z��Z�����L2U3����l�L?YV��5A+bQj �&���ܔ#\L��#�ɯ���z�g���s0�p��q%�gD�P��lWjxR~��<���m~����DI����n�`[�%c)�66���$��Oc��D;���ط�[��X=��K�6�35���q�x��XP���l}zd�� Mtb�+��>oV8a�"���^���{����_J�t���6fъ�����}�������0�6c�݌�~Q��{���PP}��Y+���00��\��ϻ갰;/��+�ٌ�=�sa �x.��(Џ���'����)9F�/��`%
0#�S����ܭ�B�-�)7����C�/JW���-�@�~��}�@���P�p�����[�������.�C��0��3N��_b/n������EN�բ��e�B�z˜+2b�����ti&�Q�����Ob߀������<����R3BL�4���8�ӭĄ��,���!-܅cgw-y�yt��3fM'B&��k�5��h/
$A��c��3���KՈs���
{��3�W���տW�~6e'�N��W�����VBs4�3'�"���eÄ9��h��ZK�'��"�IO�j�`���7����.RĽ�6)H*�[�ٲ�"W��r��\�3��]�8��
T.�b�ªQK� [q7�����vF�0�/�5-�jdl��"n �i*���� aP2�s���)S�d�x�Z�Ң��N7��!*}'�_�� >�GYwJ��X��6 �g�u�u����|RW:1p�ש��Ȳ���p�'����q�Om|(|�>���Ӆ��h_��,Nԛ���ێ����'/ͺ'�"=�I!c���� 8��j�[8ǫj�= ��)��<P3P�$q�I��(mX�"�!<1�w�Г�\�+,������K�.Ah��&q�JcZ���mY�s#�8�r��bU\�g5C�Q2��&agz�$�i�aI�I^��=6����!u�M���qs�;������I_M�Syo.�j`~�:�P�]�u��F�ѩ��rVć�.yE���;2�w�0�v? h�L����0c�U���d�V�7�п'��Q���a�J-�?��u<(���>�mMF����3���>Ch3l�MF�^���!]G�#��)�o_�%�ڸ�G}y���cU�/�M��jtn�g#�O���������>X�7��&�+�6 �K[��������EW��[�M�[�Zv�t;sgmQ	
�'�z4o���[���v�aJ/�]�y$\@~�Ԡ��ix�j�����C���E�訡�����>QC�}j#���éDӚ���5j�����|��z�V<��ՒPx.7��Cn�7b�L_D��-KXKg��ئ)}).��������{����/hzb=�l-T�f�2����ę�u�#L.ߧ��0�z6�p��C�;��hi��rn�-y��i:4�&u3m�KRk�-�0Ag�=\� ���v��H�j6*L�D�����5m��ڜ<��G�M&H7gZ�T�V�F��'�P�ۑ��Q�s�ۙH��7����<M|K�hss�!�a�:r|���ǥ���U(�O�
�@OF�F���fHJ��1*&u1����|;���Q^a��Ѝ�^we���-$�ʧ���O���<M�)�M������FP�y
X�i��E�<�g�=�����	�<�ˣ�m����W��3)��"�ŻNśg���s���j�-!+�,�D��G���*|�?��S�R�v���gźV��ȫ8��\�\�}������ A�$��N%R��v�d��Iv�ǽj�����?NX4c�,d~�ݚח�t\{Р�Ma�7z�'��A�"��cS�~�N#��ݤr�L-�o�lp���:�z��9�7��諀f�T��~eJ}������<�~D���� J��d����Be���3�7������k��¬T�>�p��E��;��KѮ��"����+x����S�4����ϡ��/:CG�­v"
��0Nsn����5���,�n;����m,�_<W���4/�[��Hi�"�8OZI'~������!�=#��T`5'�R�w�j�h����)����h֘g!��Łc�ի��>�{�=�kL�3�p�t�����k�1��4����P�R�*��VodG�"8d�������1>KK6-"h$��9�ƭB�w�_���Ә��������G*�1��C��Q�*ʏZ$����#��$lhDZ��Z�lm�U ��T=4 @0�Er6͉�h�R&��Y��*EY7�KɆy�����e W���H�x{`������E��o�X��ئ&hfW1TMƀ�O���`���G��Ⲕ����%=a�ZJ��l;�ЎNd���!��\�� �p��Qu��zz�_Ħ0�i^MP�O /Ynx�L�6���s������Zio�.C�7s��$ͪ;��|��H(�:��ɾ�^�]��|�H�VVE8��q�a���ԔM�h��^��T𦙬�b>��j�Њ��gN�C$l
<��vr�<����"�OV��1[�7���N�����+���(�FR�Ap��a�(����$ }�@$$י�$;��W��O��L�c+ᦂ�r��*R����[oڛU�Oh��\��ddS2���
[J2ZO�ӕ8�F�*� �af��EJ��o#��d�A�1,�T)u�eG�i�
y�U`/ǣ�k�X��ic|�aO���@��9,ws�wuN�*i'�q�h��o�V��?��*�J��<e��9��'<�?�fE�*|���Mo� ��44%ҹT�� ��ןD�?f���>k��8�����PL�\��U_dJI����tҢQ���+I�aᗡ��/�� 5G��K�}�����2ņ�²��Z��!�tB?�1��Ԅ2�OeK6f���޲T����w*]��_	ݓ�8��)����a�أ�<��f���t!I ��2O�e:�8�Ya~ɣ[�"|n����� �����T:�JT����>��,�-KZ�U���m�e�Y�|ޔYe�U����tg���eaS����*51�Ԁ�D�ϐ	}K���`69g�"������Hӄ�*�Hnٝ�Wh�s�K�N���H��n�L�up�i��|zR�uG���h<@O�YݥT�H�Џ�XV�l9�2
�=���3�/�s:�0��f�ߗ7*<����w�E��M0E�Q�`La�J*�I�,�����oD������sQ���h	���J����N�/J<����_`܏®�x�X�0ؤ�"����� Ē�	j
p�����jN�B��� :~0e���c�1,TQb(C�V��w���Fw���3�j,�ۆ�$���! A��h^�b�N;�y�_��;�=K���q�`R�k�m�a�n�,b%�8��g��&9g���#����f&� hT�<������	��X������`��<*��9"��9�}����E��$b�C"MC�4 ��I���^�^�D<�{�d�"�-�~d���J���w���.��9Lhf���aM���%�!�8�x$��)+R���J�ƕ���!���Q�m�~���$P�U*�3I�meN�B��Q���֬�%5���[�H��Rx����1Q���T�n�ǺPo�yqץ^�4�I���B�y��T{�zw�,�<�L�:+ Q��|@���t~��э�}Xi�'8�̛&��(a)Wb��G!!�4<��k�!�s��#.�M�G��fmEշA��y�B��C��*;�}�'�ؑ �Dci�wNlX��W�ʼ��HtD���������4-���.73��;�$h8#�F�.�εZ7՗N�!~.�\�.1w���r�f'{Y�,�;�o��o����{	�۱�pˮ�j,�����4Z�?�+|M��譓}���(c� 8�O\Ƀ���=V:2�mj�\��B�8@Q��y��Ҭ��D����AKU3�u��xjZ�����}���ڇY5ط+��e�l�L���q��[���Kg��.0��q��`��a�����svT:�s�H6�{�*�Y����F�kШ¯q�M���fH��|�&��Z�\E/���D �(��nv�Iy��� Yt�\ �#Z�}=S���Q�6��vm=t�jD����tʁ��w��  _��N�[ճ"�왯D�Ĩ'��q_�7,jLL��f�a"n%8�1 ��<4��8��F���<q�8�2d7$mи3�e�L}zE���@[Kg�l�w��TX�2��}@B
O]\+
{���^dN��N��U.�D��YvlДR��� I���:*5�=�v��4�Ώc�mJ1Q����fFy��)�([�2N/��unoR�s9�eH����]^�{���\4w�Y��6��������^s�iG&�²��ӫJ~ӂ��,�dwfk�,��\#�w���k|b��~�v�w�,�7��e�ͺs�9%Z����mH����� ��ш.i/�^~���~q
X��pѦ��e��(��x���xz`��1πf�!��"�_�y�U�F����29\DbK�v�V�M�L��<�#ݑ�)���ב+�?r��߃���̶�K+rULgT�t�_t�G�.��u�s�"¼�f�/z �ݐ�^e#���	�n�oNO�o��d����4Z�mV�C��<��N�����!5_V�wnN��n-{9xʚ)��ZIfĉ�;� �O!�_2yWv���Ǯd��Ց:�K@�ꬦ�K+��',�X�|c.,�ƙ܇��d[�]<ŝ8�^)}p	�l��U���"�K�u��L��I�4�E+Ƅ,�G�������J������oO�a�C�g+v��V{�(�-o3��{���\�P���������Q�:�<O�������'�P���iՖ׊ف�*���t�<Ц���r�ȴY���g�t���Qr87���R%��w'�z����2�;�N0��%0����=�E=뻏.T`Ξ�z8 ƚ5�=�,݊�i�g���^~ht6CkG�vI�����Vv���j;J��Z�#8g��W_p�0Ƀ����<(���&�0w�	$��u�ǚ}̉��g�a��?n ވ�&�j~��y�K��+�"�#�L���8K�
e���J��/:
G�2�3uG���yc����A#��<E6���O7����3Q�fC[� 4 ߯J�ԯX�0�J���-�|�6��Z��Գ�"f�V��%[um�u��p��㇠T:�V�P�tx;?<�(���\S&�E�=ܦt'�P(N,x��H>�K�7�Զ�%�G"v\�)X�]�Q��@lk5�/M��|xU��ݏ�$��DO��2�t�H�}�e��'�dm�or0X�*�<\�ipҼ`��}Hc���6�+� ��˭c$;>ח4��6�����f�J�Dl�"�W�N2-i^;L���9���-�z=�,DS>p��T^�a3��=j;m�:m�>t#Jog[�Y�!A�������h����|��<�-�D3Y�󄀝d!���l<�'J��a��U�A6��8�Ö���5�/��!�9Q2?*j�����	S�� i���cΰ����� ��=�V��x}�%F�C?7���7C5f*�˞�-�Q�֑�p`�B'9�w/��1!}��XV�����;5\�?Z%���K�.�q�	�*gDM?�<��}nL�5r0�o5���0��o��]��_�u���À��G�����e�H��#�-�qe���-���Q�S6�����m�Xܟ���J���I�2�����jm���k��b��F+����5Ut*���2���p���*�����agO%/4Ж�轓)oc��H��OZ�@�_|E�˕S�S���*��K �I�{��ʝq�<w�+�2R���r��+<��1�AP��h�G�Q�I8��?��*������qHC���N��#���]br3	)=J��k!ت�p��Og-�{�x����1��/DH�6fr�5���]�e|��O\��g�8�7���Lc�Xl�_��5#~=Y^d�!��N�z`Q�ˆS~���=�j�&�wO$;�:z%�HU<�Tک�ǸeN5�G���1��/N)�� �VZu��C�)�1�,��n]E�*؛�=K��K�;;�n���8je�s,�uƲc�]�1�qj�6
v�p��=B�����������v��ҵ�/
y�����D �ّ̉|H�'qL<�7�(����B��8�L��l�M[��c�E��jۻ�]�L�n
Y�<g:�g��n*orq}��p�]�6�O���H�s&�@Q�/�Nw�S� dώ$���sA�QP�:��&;�4�0��H
B�y�be�n�?q.�]�g^7��X�ż���w�!�͖�Ν'�K�H�՗�^����F`
���/���@&c.��{�M4/k�^>�l'M���W:ߠ#|�a��Э>��Rz�_YI��|хIP����'b{/�"{og�{�{ߴ�yy�É�f`�
0�|����
%_���g=�����=(�'!�O�W�E�|T���gz�YY�֝5c�~M�MV�ؽ^L�5�c�gT�kM�Z5 &I�2�������4�'�0�_����Q#�H�D����K��B��Sml���k��bP�'����n��"H8-����(���Қ�;��E�ɰ���QА��$�Nl&Tڗ�W�|���͖'.�����J��[0#�dA�W�c�܎��0Ļ-�Qs����d3`��f{/����*��{�	� z1Ǽ �����(jkr��;y}�5�Xra/��q_g]����W]V�9J�� �Y1,נ��-q:�D���z�'H�yg7�rEʐ+b���c�0e9���Q����~!/�J�����a��:�1�_��O���*�ؕ�Ƿ��V�KNjƴW���Ø7���R�?�l���`�T��4��������s�J|ؔ�ţ�+�¬S\N6��:�v�;i�?�)\}�h�(��@;�y=f&`0`.�B����(]���Ƴ!�w��^�2��xG]^��6�8ٰ�.fl�]@	T�+|�����^F�&�; o��[eT�A�d�`oc�/8�'
s����p�������N���� v�Y��!��Y�R�u�y��3�M���}W�� s�ii\����ID�b Ğ�.f���Q/g̓�� ���j]xUj��;!����̌D�6����\u�Z��tldI
y j (XH�ㆤY&,D:���WI�HB�b�F����1翑wp�>p<�M�j��\�A��.P������=g�x�u1�������.�+W���+Wx�/�=�P�4�Q�S�Sr���>^��r��qSl �?����0�3�Rc�z���}�S��%�J���r��8�3�$.����	���y��5�♷��/��n���'p'vM
%���;Sr���3��]��@q�� ��¹D�u��}
k�b���?
>���W\�FO~e���P��Ji_~*8�+6�[���Ӳ8�_E9��n����&�f#�U���gz�.m��;/k�(���5�f,:x锛lX�s ��'SLƣiۭ�O�	 G5k�=����0���|�/z�u��;"s���x~���ã⍲�>f�����d�� 7�t
��U��n�U� ��|�Og�1��X}��R10�ܴ�rg�m����]���fc���� ����4�W1��j�����I�j���.�Y�(��iT��1v�3ũ/��'%Qh�E�W�T��~+�A��Ci������ �Z��%6�y�m�/)���?�EzEu�&/�U����P֣���H#���3�(���Oc}'� 9��i'sB�P��}��>��b)l���F��Uhj��c�	�~�m�UN��T����[�ZX�0�D���ⶡr�WR 9��u�-�^exni����ҧ('�(`����y<ـ݄\3i�$~E=�⩬�����<#L��c�M���b <s��A�8ĩ��}�HV &�κ�������s8¹���&x	��w5�6�J�4Cv���9�Q����`J��F���Xu��V8�<w�$�����Y��+切Cܞ��}����\�լ\��( ;/�t��PA�����x�o���bFt��_�$���[}�g���0Z��{��߆>8���]�J��y�Ÿ��i`�Ƀ�XL	-��_k��I��3Uwl]�����e煺�����Q�`<�j���g���u1'ʅ� B�(	2-U��s���Q�c$(/�� �Ũ��&��[h6�x��w�!�k��u#$�4����@uG�3�,�,F����g��#�����SM�Nk=>��UR}pW%����IC�򡀵�D�9�o#<�S���G�=t)CiC`co�P�(��,�&YϚ��C����H~�`W`���=��̖���'��/���mҞi�i���MYbCF0����­ں�>G��]���x$I@ u��(;K����t�&�,�_sWb�~����Q��.Ϩ�N�2N���1��y�^����G�9��k�~+� of1�5.V��Pٗ��*i�^)gdm��&�����;��9�H>5GF�o�̔� �׊��SMމJ�Pƻf4��P���9P�����8/�����p@;;\�3ަ� xi�,�:�0��4�2lt&#u��I�����*���}�J�Xp��@��� G�2TCl���M�Ϛ���H��銏K�ss*�����'��#�$��܄���\�(j/Y
.gWO�LM����~FG!��x��V��Q��ryBj�!��2����B��ҩLB�)�Ғ�6�̧m�{�a��5x���1hYS7���&�pSV#��;��#���0[���K8�kP��r�*��U�"��l��2�.�/�s2����*u�N��Cَ�)J̓hv�:�5A���K����4u姓L�Z�xH��Bh[��7�\�6�	�{$?к��}��I_�w��c4�ԫ�[������|8{3�Z����g�go��}�f�{�tl�A+����|�M zcǣ�BU��n�QA]�B)I.O�\b]I��4�#A�~a��xE�=qbT� ���)��Bz6��l9N��}���� �������Ҡ���q=8L#��~f��v`T�.���A��K�(�R %�|�
u)�@v�4UgAGbT��-9�R�	���7�#J`�	�:h�gd���U�3/H���7�{�;�h����oY�B�`�k�����v!�3���;�{I�
�b�wL�����Q6~篸N�?�(�V�I@X�2u�z�øn�JXZ��3le�Ң_4ݗ+��Β5F����i0@�A�c4cR7�G�4L���	\���u�o�a �yrf_~+�"�$���/��
�ԫ��]���CC������l	�-�8�V��m'���X�&Kӫt���[�"2�7�
��I�N+��V<@�V%^�8k����
��k��R���t;�>�����0�"?L�:�c����Y�#}:��邽�\����v���Ϩ
Cg�}�@����g�����G⧵�mٜ	I���9KF�`ۅ�{�y�4}��>��xG����������.։`EkO��$��6˥��Í��^���2Wz�<��"f0����Prle7ۘЩ�{���D�{��_�����Y�������2l+~�#?;Z�!Fy�ƞ��O:�L���&��Z��P}��C܏���
��{ʃ:B2(Ϣ$lA,� 4u���u�9�++�L��O���(���G>���B��>�:!���06k_��J�b�P6���h͕fc�����i%d�%xʗ�na��@2!��3M�yX�;vEȿ���آ&˿��J���L��n|E6:�Z���v׺�fψKm��@�(@V'�*ѡ�N� Kq�|(�)�����gT�<�,��Vp��_��#|�� �"N#)���<`��N�;S�<	���@Wq��v�I1��Zeri��v�"|�DcZ�w�i��#H�����\��[g�˼�����6�<_6��۔Ę��I$n	�d�N�BN{iԬ�A��\��`6�2�U#����GN�[�
�a0e�K�$����J;�Pw `���KfK �'���	~��>����@n�Q��E�Sk�MT\h���M�x�����G�$�E���Z2���Mq���d���@V�=��
Huc�MX~��n5e��h�¿J*���=5�)]( }S�ǔ���#DD�$pE�0��P5h&��7y�Mx,�Z*Fy�Xć���sf<ڑ^S�/�ZAm�a�=a��"B�+\4�FXl������(ϋ�06= ��&3 ���ڵ�h��sM+�X$���d	==��|yK=	$
핖�,�8RR�u�w�K���7 �lθ;���e'��(�^.Ӵy
z_g�ƣ{��}��*qܟ��5a)/_�W����
/Ɣi��Ss]���_����p�uo%�w}�F��q]Ҙ��-	s�Rm���:5]�%��3��F!`�����T��#!�aY��Nd�9��BZ�����s��)���ɪ�P����d�Uz����v�J��By,'M�6(09$�-��J$A��SFh�0i�����{J�O ,��F���q�@P����bb��8���h�Ġ��v7X]n��q6����D�>�l�C�С�PE��l��Ǵ�JC�[�򹱶��x�r^c���l��x\�\�(0kh(��$�y�.پ)���ø��_B'�" 0�*���R֧����7��J`�0r����$#�	QZ�%�Y���	����`�Cq�6��ǖmcqͤÃGǪ%p����ȩ�M�D����F��V�l8������ePا@��|~���s���"M����ݟN���2A��S��!ڟ�ms2�gw�^zkyb�E���������y�v��"v�5���c���߬逼y�~Ÿ���O��r���l��1����KkJ>�>Lv ��������6��`Ni��ס%�����Z���7Vkd)nW�ͱ��B
|�� t������#��f$�:�eLZmE��Z�Z�zC�*:M���%]�Wī|�Z���W�>ֿ�U�|j�`T�e�|ً#����o�`�ؗ�c���u��N#�yz���*�
ˈ:Ě�>�{����o��*'ɔ����ɪN.����T���)�w����Ն�s2A�N7M�n����t�C ��'���������f�,�=��rW���%]��YK��Q�G�E�}����
ܘ��z[Ո�E�eB@�Z�B���ԋ�u��qʗ�k`͊7>z�2�\/�rd���;�L��[�koG"*LP�jA?���Z�!���E:)��?nD����V2t?ƀ��KI�E�t�2�8��ᯏ7�R׺R<i9=�{g���� s�U%�ϟ~U��֎p4hŗz�Gxv��"�d�[b6�+8C��u з@4*ɝ*��Q�g�3@�"��(�1k�r+�4g>����i=[�{3��\���+Cr�ױL��@�F��Jٝ���8�D��4�C�B�K�4ϺD#��Ζl�|�G��t	��>�/'����ݽO��(��wK�R)��C�J@���<��Ac��W̓�(���V�$@������mG.a~7��3V�1`n�'05�a�PPM��T*��8��uǪ񠶬�x6��
k~���f�o�:�Ay'T��d�߁�9����u#��)6��#5H�E+��=��%8�D踤�|�c�L��9 M�4Mv vͩ��Ы�J4��+��V��=c����:��rSҽ51�ԂqF"���I�7g1+�)�y�1�'�k�i=|�)�Q3�����D�3A!�~j�fz����#.�Y]BcA+.�+�Z����#E(gM<�n�ND�$$&꽂`���-j��K�M���	��Ӈ�4wބc���6uOhv�[���L�Ҍ/���@���\�(�1�üW6oa<r�{�`��X�X�u��%�"�FM����
�nKT~��>B�ݎ�q+���#���[:V��f�:J����o��$J�N�+n�M�l
@���fv���!]T"��W����@�$���C����\��L��n�P������ϐ'�:u�'��-Bq�@]_u]Iһv�����w7u�<�$���|�D�_9ж(O� 9�G%�;����+&�RL���+���&e1hRMM��맄z�E�E��m�����n�'�eV��E�Ɠ?�����H�I�Pme�<M���`����~-�Z�m��@7�E��Eg�%N���T�y���Q�Ä�_[+��Td��6�	�

9|��gy4�=���<�uV�5�8zi��!�UX���f��	`���[ �$�`�6�NN�I��>��$϶~G)ZD6�&��'%�*-x�R���{+FN�il%���b:{��l6��ٻ�s*�P��UbZEڃe2i��rp���zVX�f���jz �F�y���B���]��w�B
@C`��$m�,a�帅���O�7��2�؞X��1w&h�?/�^;�D��]T{I�~��	�L�	K�����S�=�@q��Kg��(��^RK��w�$�;�<C�@uv�X��V�u*z#�q�^�y�����=�9��5�̒� ]?rG�zUD���;��u��j��IM1!]�:�Z��:�iV��E��ͮ��ր�_.[7��ӍiGNB�#������$��bm"�*�l��܂R{Vf���Ň}V��'�lM��/�&�A5�8�>�!խ/Թ�9P"��k��z��Nw�>O=�[��o�9��E�6���Lz���|o[��N��
g�V�i�^/'V�Hzh�?�C�.a����G��,y$���F�L�r�!���{�=G5��/J�#դ6�����$ۋ`�������(��/�%ÄC�$��85,���<���=�V|�`�������59��p,�����`ȲIxX&��Q��u�N>�D���ur�E>�h7{��0�r��sUBO�׫ˍ�ڠ�}�y�ū��1:6�#�fS�䅒�>����U̚^�0_I�f���f������!ೳA��D��=�������I��� Z�;r�~1����$5�R�+]M\�.��/�e�&��7>��Z��a����%��\q�?�`'����R\��e�7<9�}\��7�<ꆵ#���+	i�r�����o�1�Js�$�/����^���QV��각Ⱦs�p�J��"ϸ�o�/�%}��T%h�:ΙxVh��O�H�`�b�7��E��޶���	�(�ޙ�(3���m3~Gx�� _���4r n,j���sZ��JB�MX"��?z�t��eXmİ��4�R#��3HX����qÜ9sLDɢ&�P�~x��{HoJnK�*�W�o':������g`N�W;
K�8��$,�(�xw�]�$m]w�����YAY�j�i�1�zr�O:'i=jfl�-���# <V5C��lV���
��k��F�C��u�yB�.T��`�.,���:�����я4�aVW��Éq�>������7)*w��h *Y$�n0��h�O���%A	�z|�H�,��e�j1�Ȓ��������Ks�ƿEDYS�;��c��jW�V���_�L!HC��L%0�h4�m�P�zn�?��iFz�>���fʂ�Z�C���w�\r�&�.�<D���,�G�$���	k|�.�/��ә��΃���,��w �S:,��0��N�>��Bx���a�}&�gz��De`?[ޙ�$�x�w�Z<��E�GO!��AIu�Q���[�Yth\?��躷�ZA]3𮁙g�7*!�}�nK�L	@R{��|���,@�	��ԫ���L�B�t���J��e�l�r���@���V�� $��������^^ՙ�+�TU�S�1��lh,m��+1F:R�뻿�����F�`:������9-X���c ��9�x�bn:�4E�½A��7m�BQ�B��n���$ܮ���t(��ݐ��?�'� C�<�� ݡ�`��gw�ѽ&�S�<��ɺ��V!Q�h�+7{�F+`\:|po�����ȃ��bt��s�U@�f�tk���T�!���Ӻ�8���g�!������aI�%�ۧ4ڏU��P�\0w1-����A���a��
��߽J���U�h�n�N�.�1��$>�d��ʻD��;$h�(��W��%H���ِ�6���0�`8�u��wz����K`\Eӂ i�#WG��f��%�.�ܺ���w���:���T�r5:��"Z	��U��{��@-{GE�!�sv������a�G;�OϚ5;��O��j@��1���^��wZUPRPd���ꔚ��n�t��3U����bu	$�1Q�}Elx2M[Zx�֔�RP
\�
f���B�1ǭ�a�|(-�37���ȸf������[}�h�plA�4����b�=��*O���2�Y�ù9z��-��FD�e��+!��aU?A��!ZPvP��ޥ)�L�ks��r�E���х �Ci��@''���cQ(����|r'ɼ�K3����[�P.�3�g��$Ske�|�l��\#����L����z^=$�3��8p���Ġ�-ܧ�~����l�f��Oh!�0���E��P�V� 
��7�3��H�4tF��{��e��y��"��_O��Oo��WS
'����k�s��}�~ J���)�U�.�C<!�+�[�{ ��ܦ�k��n�7�wL�_������ ��.OE`P_���5��8�SH{���?����� '��"j�l�ݴ�1,����񔏠/�&��F�'�s������B�?�x�xKW��W���D�tp;��ouЉ����CnA]�v\n^#��\?��Ϛ�]g�sx���ʏx���8�����/�<X�\��Q��6bY��(��K�pPӓ24}�k6�A0D=��ݾ�;���s��Y�����9�E5\��pۣt�^��a�Lʇ�U�v��;J-�Q��r�0D�3b�;�L�E�u�_ң��;|>�"�cg�ҧ�I�g�մ-ik��8�l�u����M2��;n���9�M�# �P�0� �{/�&��ɉP27�1j$:����ވ��zKm��+4�-�D�Ikڴ^����x�R0���`�L��q�٤A��toƉq�k�ŧ2�#s�Q�,,�H�6l��ݮO*���C��Q�aɍ�|��O�F���\�)���	�Ô���������Q��F�>H��������0���j���\l��DE��-U�qL�w�Wˏ�%�d.4F��_�oY�f�Vf�q��?�"���d�k3��U�ßpL�<�	��Y�_>�^�η�ޓ�t*wp<�g+��aA*��u�ml��"��V�+���5Nl�(��Mdz�p����u�0c=���^�LpVlGSi0�F�/\O��GV�h<eC��)e�0���,��F�6=�[D����1=Cw'�s��9Jb\�����X�z��X�^����鍎��WTtn���ɬaTb����p#uADRZ��9�۔����x�����*�sD�Se݉���j�M�3�����)>�����q�@s���a�2� ֔��dBRg���3��OJ��#[�I\�^C��r���քM�̣2�H��
�=�N�W"G�:�D�2Q����?�93�G
:,�感B�Q��g�t���4Bx#��;���3d��ŐE+z��e�c�0 r*�EV���_��g����q%h����M� G�Ҍ{�ѪV!�>�΄wW��1�]��ز�	� ��Qy��M�!���}B¼V�������^���R���x�L�����
�?wF�6,Ą�E|�!�[�;[���~�������i��]�<��OR6p�oT�&�<@�Ÿ��i�p�d��!�ƃ#���:?��6�G(�&���p�0��������I�L�ޝ|��~���z�3�qEPv�hţSǘ.u��e�I���1ѭ,R,�L���^ʌ�R��'^�lέY�Xc���e�h�nx�s#�+����:%��G2��y�P��L��ͅ�q"8�︆�z ��f�L#"L����o�y�ҨtF����)[Q����DZ���d�G���3�E¶���\����g��������Ή�
Ŀ�J2�9�k�F�F&G��R��C@�j)k=�N��7����T6x��2?	ؖ�s�U̔�>�4��`{woe��e�&$}R�:�S����G�QJ�������̮�k�NJ�NI�=�w;L�!"����}�@O�wH�ƌF����Y����Xu��������w�"�l�H̪->�hl���Mh��>����r��m�+����&�2�*��O�Sdh����H9pX)=�����]����,ě%l�Gg5��e�7#	���6�k�g;���'��2���;�"1��Ί�]\p�/Φ�A񁀲�JQ{�=�Ǻ`�8j��;�Qm�7���y�N�ղ���U������X�DT� 1g������x=P٢�1v��uCC�R!Y���*�C��;�\rI���3U�Gµ��>���VCh����z1瓼#W-&K}5m� ����:D 4���f�Ǔ����TB��⮿փ�UY���� R�"@j�]��?�D�P�\�WGz?�}h�%�.BZ�x��ٻ�|��]�&�&�r��$��Do��c�����D���G<�=3�{�'�?IT���l���E�M���/=`:�Hltm����X
.�>I� ��|�:c��1^S=���i2�`rPG!����L�`�O� �1C�G�_��{R�7?�e}�dƠ�=�J~���ˑ!��;����-FbX��3j�U�Jj�%���Z��z�@���W�6F��M��\��#�clԵ2�����D��b	f���"����_�q����t}��ec��2[��Ӻ�=��Y�ͼ��/~��u��k:��IZ����8.A�ޤ�E�cH���0����B%EX7<!1������Ϭ]��{wt\]x��Ձ��HRg�R\�
&��NgGtP��d�9\� M��|Wi���~��S{e�e	���YSU�7�`w� �\E�kܙnV��C�D&X7"�!���6�Ǜ�L*l�P{JX��H�������G'�6ʐ&���[2}��C_����#d�O���2D�vbѣjf=ʵ�S�um-��cP*&*I����.C������G���g<��N�!S�rzL)��"m�DV�=���}gM�>�#���>���[�2�q�#����X�lm"�~�W��U�;m�;��W��ﰩ�J߸�qi݃��Y3�z7���@�Ǫ����AR���Y�s1����{��TP�}���9ch�I��:D`���[�h{a_]�Lr����.%b�B��wiέ�ު˄xZ!%���O�ُ7r���֬ŞD�����F�CM���1�B�ۏ/5q_����ľ.��<7�#�bW̮����e��m�C]���>h���`��=q���F����v����<`l�vq����x#4�pN�?g��k���L�އj�]�R���/�?XS���f>��9��	��r:q`xRA��/�z�b�U�,��6�˫m���w����O�`�gkywN�#���wl��_����~>��MsR���.���32��!�%/��o��:�\:�� s!�����4j�{Φݧ_�!	ږ�y�T�1�_7�G�c1u�VL�k�Q`��iQ ��5�����ޗw�:��:ϲn0-�ρ�L����\�O�\<�ܾ�_��;�t19-��`�k6E��%�M�&SE垨J�����f��wk�޳���A�;�� ��=L��=E?%��,v�nk�Mه+A˃<go&q�����+�'�Z�crTBRR݁����bt3��z�jYlzZ#����F��,�P����P�o].M.7_�e[B[���p��<�и��̑B���<{t��%VSӅ�`���XMP�pU�����(� ���%���@�H%�z4i��\;����Eg
��Þ�O4������z ٟ��બv�� �R��iug�Vw�{`9��d��Zu
ˇ���v���A�[���$|Ѐ�}�h��xg��?�D���1�HY+o��J.�m��N��س�I����= ���2:]K�<�AO߀�!)d� �Y }��_��do�ns��W9��\`]/RL����%�0�P�T���!��l딾Nϙt��Ʈ*2�������p�k���hUT�,���Z��x�E���?�l˫Qc���hkEE����m�(�QI7�qg��8�^��K�h�����}<�2��v�/��D�UV����K�334�m\���D8XQ������4&�����x�(K% N�W� ���<�h'�X��rD
6��ud��
�Yye�X�/��4�0}4��x㎗��As��xA�4`�z�|���47���=���Lr�֛�B�ǎK	�3JN����Q�A�~. ���&԰��a��cN$���QP�L6���+���{��s5_�b���-jz�^�쑳��s��l}hn��:���S$�ƗuHR��)�g���s(�������q�;���=5�s;�_�|��5G���������,��$Yk #fk-�����bȆ�T�oy�eX]q�]��n5�{���9Y�p��ѯt����2��+�� �m�6s	��*=��ØW��d�luݍM�ݝ�/��|7@��C�����"��-�b�E���Q�yؿ�i���#�&�DM~��L�t���`�LdTTxCF¤��˩hʺ��D�%UQ+�JNMn�a��-�ׅ�o�B)@t�1c�B/0O!�3¶�Esq���C�'*y{-����G�̘�A�7qo<����ѓ3�V��{�^�Q�+8rX`���3T���Ո���崴��(JԎ�Oz'�[�aFrQ~��i!�$.��%��E��i]�Ie'��`� z���t��0��'҆�p�x�pщ9 *0���9�f�/mV��HSI�.ַc��^��~px<�(�}`�i��ÝFnk*>ؙ�;��e�|���A�:�����������C�l�P
��S;����p4���/���h�KT�ڈ����kp�q�	^4rn�w���|�Y*��R����x�4 �k����.n�A8x����Or���_�^�b�U�F+���:h���ǌsq���N(��.����:��]$8�{��)"vqB���BjёӍ@iY�9�Q=[g��4�Y�5�m�l�ȅӄ��R�2�Z�)�d�IuK����X��*�'���je���*#�j(z��]r���rݏ�h��~�v*s˭b}��({�Nޥ�X�mo+o!5�'ڃ�ѣ�^>�����YՏ�t��2M�ױ3["Z�M����j��]AR��q)B5w�w@�O����.�e�b��ۘ5��_˱=)\8S?�~�][���~�c봳�}-"XJ�$�J��`^��h����<�(4��gIe
��b�ҙ�ƈ�^�9t0���~.�RS����|�
J%j3��倧�C��-�Qߌ��Z��]A�q�\z36���Ǟ���)����c�3��ɹ�\tn����o������?���E,�N�̀_�}����eXh�v4j��Ÿ`k��7�Ⱦz�>3:W����[���D�t�oN�R���E�(��xt�� 
a������X�49B�C�5�,"�Ó�)��ۏ<�_�gh=��G�����3c��
���k��z��/r�:Ψ1~�$�1�hH�Kh�@s ]#z\�G(=��n��l��NFeE�_ӣ���mc�/b]�������U$R�Y�M«}�"MTl�,@�9z�����vד�|�#���C8/��,�=�7��	��V��V�}����t	r�}'�&9#�\���i�#zԆ��ZX�/�(��Tml��t[	t�pA�L�S~K�s�A��PRB�5e��f@���%GP������JVPl=�����)Aj������e��r�wr&��:Z�|9��vO7����X�}^8K��v�0������,���G=�ex�i*�5�Ur�)(����+��v涪¢���]�����	�Z�Ʉ�{a[oZ��4��"�3I4�]�P�u&��,+<(5'�>�M�'w�h(F�D�K�a�E�����A�@Qp���������QLF2u#�b�c�Z�(h�}k�G#�@��k��)��� #\��gX(��j.r��xfM�!��C��H*m٧yXݲm�!d]��)� ,�$[.?���ж���q�31ַW��}tZ���Z���V�������{�ޮ�?�~�.�#,����-�N��xλ~T>����� I��C
���Cnr"�<?�T��d��� Ȥ+@���y�z�����
۞�z�7�W_�Rb����K������>�ߵ0���T�	Ž-#�����x>"�Ln)Ay���ZC��&���j��1aLm2�Q��m�Ű��a�V�D=�8_�

t~H�۞��*zb�Ԫ^�B��e�������n!藻Y��ԅ���99٘i��Z{�yE�I{�`	�Ƨ�m�A���m�x���kP�/f7-jCܭ^]�i��_�nw�L���vi� X/���( ���Q4+��	=��g��9��Қ��������h_���/�r��#��,�sP���bO�d�=�*�J�r~kc�h.WY�}9g��9���[���On#�r�@4��ȯ���P����>���е�����=�������gŨ�qv�d���_���O��kqs�{��˦X�'F�0�|~A��ǹl1���rV�QW��D�q�[�]UW�5�cy�A�
�%�GBC�E7�����/�E��!�u�Cnŋۃ,˵L�q���l�d����w��;��DG`��l6/m��B����1���Qs�IGC��@�GI
��`���As�_}�8�0~3����56I:��RB�ߘ��᡻6��(6ϱ[���}���g󙆞�HB{t���Zk0��_ĒB�� NDf��|��@F���%L�R�`��+��^GC£yN����	/W�c�dQ0BPs�a������.�]��fF*C:�P�yZV7��l܀����0_�K�M���V����=�ג˒Q�e��5tRud���}<~���d���bi������al�X	O���j��}�\?3S��j8_#��d��g\�1��0S�iP���ą]�;�bW���b��2g�
�l�:dʙ�o��J ϱ��N~�O����Q��F�[~('>y�� �3qZ����{z-(����g��u�.����e�#�}���ܕ��-' N.h2�k��H
+��L��4��mq����aX���K8=��S�y�� l�-���qG��r�+�/v���Y�Ep%<h`͖�÷%�;��>�V�Ym��-K0���$�e�.DB]��J	��"��]2�2�p���猠%w��6Bڵ���B`߶���5�&{�Ni��b|;ܜ�4�W(ScG��)�D�*k�P��1㻆���z�si�A	�Sp��É��3�f�������HV���V$��9�P��J`oQ�׏JZ�:���*��*���i�������E���)�����-�9����>Ϥ;or���y*HW6����ꐗ��)�[akD�eO%3�]����*�~}a��O(����o��H�Kvd/�a�[�Ԃ��*K��P��ws�M��IKp�~>/��"�������w(ueVT�&+�0K�GO�U��ڌz��b�T�M�T~��M����g�R�Yi��jb-v���)���Z��IU���M��������@*(,)ߌ��"ϭ� zlŔ��x�5,�+���1�U(�k�B#�D�w�PF��2i/clnYRxPQ�Y1�3������v���u�ȕ)b	_��Q�f Ʋ֐(>)/g��$헇�.�e��.�4 �����le܇��K���)G�Cq�#M=���,w�v9
��c�k�1����\ߕ{�4G7_���!�E笂	XD��tG(�s	K̭"�3��\mL3�s�ᇟ���F��D��=�k�Ŷ+��,�8�Ʋ}��C@�8<T���P]2_��r�/�0P��JB������ �6����s�}�`�����ֽ�1���B�����E�� nn
�MZk�o��Ȳ4����2btR��S��93T&�S� \�l��|7�2n�^1ք6�=c�)�T�)����[��Yzi�{��zfH˫cL����oP�u��2���ɤ<c��9(O;���u�X�?_l�Ӕ��%۪�7�Υ�F:"]����B����qb��aW��i"�~kʩ�?��h4>�c�iS�IB���g�DO�D�	yMg{�?����'��'�]��-���ڎaʄ�CҸb�yv&P.��+ee��9�[Kc�l�� t�R�쭮؍�X�p�.�X�W����R�g>�q��Y2ڦt5��)qv���4�����q�:vso�V)~o;�Fg���~ٺ'�;v�('�n�	�䢯�U:�5�J~&;��Z.���_�s򹆨��
�JO��.�H`BE��X����4�+�K�+���y�ϸd��Yfa�= P}(�8q@{��S�ēe>2F]��v{�g�I��;�7�R�7�s-pNS3���c[�Z}�YQr�b��Tr(�V�o�,��"P{���V��PF�x!%�!a(�C��p{OjR��g{�˛���̜ ����c� ��<sG��@����<�Cu�F��PV�[��#�n�O���d�l#]��+oJQ$�K�
&M>0inl��Cx��vW�R� M$#~K���]�Ɉ?_�����ޔR�Ɠ<��b9�+{����2�:��hJŅen@�ݜ gr0w�O������	�E�P`��>���E��M�CY��(�"� ��x�9*��Ka����.1ήfO����W/��ہRz!����~8�|�
0�x�^�ME�߈�cE_\fh���������K5���ӑRez�(���]Ko��C���>h��}��jV�������Տ������B?ќ^���m��co�8/w�)(E�~�¢�`��񷃡R�����|��2� 7���l��R7�諡�m���W�~t�ܨ(�_�a5���C�
n؉����@$F�/;���ME�n�f"D��������EM��a�NI��ﲻSK𴼝��f,�[�s�ޞt�{j���G�R|���g�x)�G�c�� �i���]��L�E�'������*������$Z(٫�U�=64�?pg�x�H��/������G���X�CT�IG�g5���JpPE(��ik�i��/�A�$�T]�Q�S�.*22�e��; �c ���i�&%�ȩ�t�& ��{AVH /+:,�X��Ah�7zy��� e��1���/zxg���!�~"����p�����mr�FT�g5�Ӗ7��]��R:�f�˲6F%@�؂xMF�x9��x_/����d��Ĵ�{����a!�=H}`��іF����G�a[�j�G�؞B</q�E��� ���)�0fŤ�l&vWe��	�v�1)��v�s�_;&��؇H�)��[R8��?��_���������	��U-sQ'��OÚ��@�W�Qi�ލz.Og�/�<�I�:Gui����W}�&��,�aE)���xؿ(�p�3�˶i�Bݙ.��|Lw�*Jo#�S�kU�t�1��'�M
��_���0�	<���o/�@pK �b�x.6`�%���|E�n�(�����F2Wa�mǛ�k&٨�k	�_Z\�r�62|Fǡ��n�Jk���B:�
���aL�JDWm��t:!���5�1�F1��&���.�U�\VO��S1�>���+�P����Y ����=?��M R�-����"%_�/J���:� �Jj�"�e9<6��D��\L����l����z�~=��YbE��h�m^ݰ��9E(��h���������+�l[k4�!�{0�����5��U���W�}�����g<�K�ΥYz<e�|[{߅�����p��~S� �)*�-X	���5<=��Q�12�VCD`M˩��/}E�hJ�.��`�%pp7�\8"��'?IX�f�Y�7g�q�=,g��F2�ލ��C{���t��ɹ�Í:��E����*W})�Rۓ��"��u*ÓJ�h��[��8�0M@	XO��I!�5~�y%������8�5�lq�����x[q��XB8\���[+�8���|�0��w�-��p��'�Bg�"l��{�~�W�t>h��xrs��q4O�Uh��z3��tF�J�d5��-�������X�x�t<Yjσ#�[�^�:p��b�"�+F��bC�2�Dy��>N��7[�}���B�Ò�5�py�7;09��ɤ �g=!�gc~ЃU0sA& :� �Lg�J-ͩD֋gy�?�`��[� ��6��Y�.i������2���K�ŅQ�v`�����j>*�g�x�բ�"7����8S6�˶5L�8|BT���2/�f*eR�ݎ$�� D�l-�m��В�!q"�#�NWR��n��ܞ���H����v�j��N��R��cSu�Vg0R��2@�X��^��ׂ~�6����� �{�\�յ�_�TP8����6�e��)$���Fg���Y���\/�{z��Fp�����H����e��O�T5ߐ{SG:��F��Q��3��!$��	����ܫh�!��4i�
Q�sy$P-�ג���&FHZgf��	��+,� 덗�8kv��x���$O5� �0[�?Wx�{�g��-)��S��VR�y^y���Y��&bdR�q�T�2�Y�{S7��VL�@�=>ȫ�+)�f�ؽH��������UH��'�E��m��Q��7�u�J[#���~��"��j�0�V�>�yE��V+Tx���"�`]��6{@�v/
�Y^P�r���7截A��^�@���Tr/�N�r�}KZ-�<�/lE�3�_��	ӼY��_@;�\f�ˉ��g�CS�^�>��~��O�+�_���aeK� Ao����?9�1�yZ��?'P�3���]f]�ha�"��>v~�2�M� g��g�/����G��g�}e�:��7�n*��ȕ�pڰu�ئ
��o\/٧���N��*��\��Sl1������t`2�N���TK�|�������5PCWY��y��Im�־{jt���M�1#�`?�������������s�.�2�m1�;�L��>t��<�e��/� �_��@I�'-I������ �+��8GƍP�$C���d�fQn����e廄J�N�J[�w��Ր	� �&xf/Z C�`*�8��A����Ԟ�4uPS
��:)d={������G+C�	��2�4����G���ZD�Ur�o%k"�0ސG��W��j� �}B�[ȧ�<M}%�\����?�� ����q�a�B������N���u\P%�M&0�_�NNӯ,��|�zÅ65"rg��Ř|Nr�&�|��n�Nj��O���B�(��]��Z�dMeq�|�����<�P��9�rXY�î��9�w��w��Xx�ʱq����>K5���.N��#�\Ӎ79����e����O^f�un�N<��V��m%��1Ay��i:"VIo�5�N���߁:������_�KG(ꏣ ���N�����L;�sVE�e��;PY>�@*������ %Y���7��� r��8�%�(��<���f_�a�P�Y�Lc?��jk������&鈑��I�IDHUf�̀�U�=��w��D��/ \w�ȑS�$�R˛6׃��uj�wF��1F�S�?��H/ʧ�X��F�zj��o���D�$�oy=B0�i?ʨ�O���������^,���.LɅR����A�7'���\��X�H�-���n�N!����1	K���
�c4uŤ�x#�>���)]��eD���tLۑS��0�<koHs&2p�vI[7��o����@+��0&�!2������ &�S\-�ZK�ޜXÀ��1i�C���Hsi�v����zA���U�ۈ�z�l�:˺wy&)��������rL��|p\��V�#�V�2EҺR�hA���n�Ȟ ������VГ�:��QA��!o����ڏ֠/}��etq��!ux�D�$�q!�_7��V�#�u��H�6C��&��l��Z!Y�&���R�,��&	�<�S��$�T}O�oH������j!T�F�Y���K��]��%�HS��Bɝ~��kj�%Dho����G��~�	�jB�|�v�|m�w�J��Gΰ�q�����X�6�x��m�͇3O�]���KJ����:׼�=��Ήu��s�g�aF���@X^@9(ݺ���uܺ=R��EGe�v�Z4+�8O��V��&��~�����ꠋH���|�T�D ���;��he��6�`,��a�^��bCe��y�ά����M���+�H̕9�K�ju�cڸ�a�'sM�*v���Ez=	b:�(rл��c+�K}-!Hu�_���L��X��q�����.j︾�{�[��	���s�"��UP���b9��Q݄>�M�V*���VyJ����,��~��
�� z��Z���t�f�
>,�![EE�P�Mv!����K�p��sr�{щg�&�tc�^-�"�����*O& Gb�C�An~����ل ���Ho��W��-xfǔ��1	x_��.��T�Np��5,T�γ���ͩ	��#O�x�1`��Q!Y�Ϡ��B}���;��_P�'�E2*��}�þcx�i5Hm�l���S)9bPk�7��0�she'�>t��׀���2N����t*�vKO|��g�B,Q\1�F��<#|��)��m�(�{�'�_+��uHkr�b���.�g-1��3�].�����u� ��3U"�tYW]"p��R�E�) C���DRF�X����%3��]�϶q(�]�c	���h{+���N�I'w�,;�ސ�]�#n�G.c��XG�mV�o�u=�[(Δ�􂷅���=�;���2<�0eR˽$�ܿɳy`5t�FD�H�.��×���{L�(�����f--���c"s�FW�y󰀅<B�&UH;��q���gEB�P���Dx����*��>V��Lku"%�LN�]��rE�ȥ�Ϣ6�%X�S�n]~h�o�W���1%��Dۻ@�x~3i��z��kNH�t"�Ӊb��RJȩ����=%� ���)4J� �����j�z̑j��6ȩ~����l��(g����X�ȭ ��nǤk��q��D�+\(���N�p=�x���l]k�u0|0����S:��>���J�0^�G�>7���l��%��7�.��B�ZQ��ѓ�抓KO���Z�c�}��zUo�����u�.Qp��>��;�hǡ�y��?QX	�/f�,�љlͬ�c����t�N�ݳ�W������Ҋn�c�)�5�q���f��j��-��,B��N:��Z7�U���#�J�lA�����l"����Eq�r�S��_ֶ=N�Nt����z����;a��P#�R�c;�}i&�#@�����u!o
	�~�K��^��,e��$�9yi�����^�g5NX�8����tNK��Mi�H��Za��{�� [;�!����3�F>��|F��'�[��&��3���@�۲�=�>?&6�/�}��Uʹ�>u��ı����L�'�L�s$�H�YjN��t��b�x|l�mm����������!�1K�(�J��\K�l���� ���A7�*�k����O�" N x@�
����ny��XI�8��Hx7:#�FC7O�Ze�!o�[l����u>���"A��j���P �A嶟�HY����
��oz��0Uxv�Z�&�6���`�����?�}�@A��7軞�2l D��_���,�_@��6_z���^v;捅9��rF�vŷ�CC��P��qa�ב���{�� 4�_�}����֖������~�k�M��fG	匀��A5z4[�i���e,�����$Na<���P�DcYտGdK�}���(v"���%)����PgPa��ќ�ՙ��J��r_lR�v��'��,���u��V�"x�۸��@"�L�e,�)�s�0�-�ߪ��oe��?��9��W��ƾ=g$ϞCxC��}�N�/p��J��-�fSw�E��{�Nw��8�%�+�1i��%�2�{>2b�����CN�6�0vI��<SY�����_wJ��?I
l'�V7_$|�?�)��X�T���I�i�� ��0��7C[��By��N�����o�`� �@�$�})«����WU|��E��P>�,��^��|(�Y���E%�������}W���T�ICwʭ�)n�y߄�W��%a�E�" �>�j``�C7N�YC�V��|��(�mU��V��h0�����ޒ���g��6�>g�hXL�]��wg��-��7,�	7�Q(,BSmb�z�O�s���s��?>a�c5�C����}�?MN
z�-rC�
����p.�\��d�J<��f`������]�N��X`�����~k�/��-��̥�:���j�ٲZ�+7�ո�d>8�-Oa� �w��m4���l�X7¦i���mm�x��-���U	ڂP��SӠ��6s���hg�Ό�[s{}O<�>���j���q�P/�1�2N/&a�]�ﶏz��w{h)T̑��|B�kڌ��%��K{C��i�n�L����V875gq�|����YQw��}!&@��Dn��i�s ��6������1�b��9��"��}D�%�߬j�*�_h���k0���x��7F���xbd&��>�p�  ���㦝�E���Ch�Vq���.�f7�SBь�3+_�t�PB&O��T��S��12hpy�ډ�:qL�ϊI"8<�hOi'`|]�9s`n8e&WDN�^96a,�`��$O8�,��M�@U^�c8��i�L��\
��pu(HSu7sϭQF�Q�>t��>�s���O���sD�
C��؜�)�:o�0E����/z@U�]����a�ܗ
��};���5�Ӊ��M�r_oC��A
fQZ�Si�k�S�kv)z��x55����+�F�D;�)'��'�by5�,��S}H�pͦ�
G�p-�}�20���ϒ��g�0�<B6�߅�v���2��ip�7o�4>˫��I�ŗ�HW���l��2<4݃����/VN��M�3���H{uqz�;�@x �Ie��ĕ������He[�A�!}$è�7<���w�&>R�[�����э�x��9G7���j�؝���-ݏ�؁��ab�@�!ӓ��{%�����9�UH �C���^7����d���%MY���x��+�����S���~�K��);��h�-���La��(�<XE�-��Y ��;�O�t�;�K�{L�>y���樱4"ۄ�!	�E�����S5�l�Ym��D�5;�t8��7�}�|~���%Qy��#,;�^z�$���/�G�)x�p�Fζ�pnM�	.�d�ٌ{Җs6��͔ql_��N9�>����MG�4v �-��7�|���y�ǾZ��.��l�Wc+�x�rM�,ULF\ W7ܱ�7��&�Z�|x]�(��Ϸ�Io5���-H���tW��,�a�W�Lλ�h
��?�3�D�lX�{}�uE�Fʻ26���)��A��%�4�+r�C�A�q*9�a��8q�,4� 9  �]pϨ����Q�lI�*��uVH[!�^��9�����6PY,�� �(�P�9j0��|�hI�`Љm:$�Bz	ho��Zh�@��Ak�9I�lG�Gl�%����"g��FQ˭m,��'�u�u������(��p�Ȭap��JbCu�:������[�ɱg��
ns� 8?�:ϻ�ҕ�Tֱ=��0�ֆq�+ez���~�v�U9?��o~��cS�S��[q���N`��c� R੐9$:��Q�螓��3k�V}�Bg{�t/l~/%�Q��x��u�ꑷ�O��_P�s���Q'�a�\��p���ʒ�����t��ϴs�Vf}_��v��|ot�y�S��"�7$)����F;�;��z����~L&�����[3��z"y��V�8T�/�.�qLors?�kyGF�i!2#� � 6wf����p�e�ѩ����[�����t�S�CP�_�֑n����-ͺ'���]*�V�� �!��UnI;��5l�V�`4�W�R���ZLG���-a���S�z�B�)5�G�����b-��݅��� ����j`��~�1d���{�eU�@0Qt�H�Ǚy�31`H�l� V�uRk�t5^��P�R0[N�)��x��J�@k�n�����ud8n*�O��*};\|��OYM�x�;��6B���݇ª�S=��}�)ƍ(<�$c�U0�
�Ji�B�ݗ�gu�V���3���@�񂧲���!%K�\���%n�lUP��P������a��e��3���65����:0E���70N8��� *� ��:7Խ���m��6�M>GB�ll�mT}e!1+���E���d߭G|����N�rv{��Y�U����/ekE/������\̠u��1���$բu�M�VU��)Ē�a!�dC���m��r�N��喎r߾HN�I�Yd�%���ɯԷ��b�[�s����U��ѳԯ8�y���6lJ.�������zG��I/ЃW�h܎h|��̢�sl=Gtgu�)���eu��Htʋ����m����9_�|��d�r|ok�,����p0{^0}
����$������B*3�_!�8�y��՞��/q!)�2����y�?�l���O�G����P)�qm+$(�Ն��<e��Zs/ (�ڸ>c����-1���R�W{�Ь���퐆3٨���A�#�z��������!���������(�)���؜iOEg�ƍcL�Y܆,	��ڞ����w="IT��� ,3Gc��p�
r�/AK+)����j�B��HJ��93��,� �����X咒#EI��"����0����k�6�9I�Cnԑs�)uڛ�gG*
G�5�`s�B���#�ۥD�t�c<���=�-�ү��.� <�3�)ق�n8Mb�)X�pt6�M2�
�V���!8A ���S`�L���D:��*������#لb�b�\��9ߴ������S�Ib�ˊ�����o�\(�8ި��>6)��]�Ə���~�\��
+����d�L�[)�lz��E�ML2Ya�V&�AW�J�A[y�sB��){Lj��Jt"�k��Y�[΀-�Q�	�A>e��j}�8�k�I s���չN 2�������}墬KN�H��_��x�� D��3Z^\�޼��g52��~�����a�"q�����!_Lh:u��anv�Y���a9����I~�8�?M�pEc��3�D8�����[r�-��-��Rc� ��"2
��Wa��;=�� c�fY�V:*ɉ��9РZ�1��#���{�1j:�_�:��-&P��ؕa l��)=Q�"�?u���c�32j�M�S�m�4�!��Od�mȯ��	��w.�j���ßc���=f�|������	�[q�􄉔�'�/[a�b h����Ӟ`Ò�tq��־�K.Jp��BXl@8]�񌤎��O���%Z�X�3��?�j ��sp���%���L��"l;h��j2���ؾa�m�lz���̆΀�
��)5[�f�B��z�DrWU�2W����5A��T4��@�(���0P��e��E��ux�&�ȃ��Q��?c��b���m�F��"��G�Vm$�GY8��)���X����'."B%�����6~��Ac�F���&��YՀ�I�-������/T�2�G�������H��?��,-�ET����'��$��c�D��ll���'Ȯ_Ne/��-B�����N���kd�{���H=����wU�78�ө|ᬿ]�)��da������])����]�]̩r�d�b�&t�~���L�GI�+b�-�5
F�mH_��|2E?��|�KM	��P��X�Y$컛�l�q��ә�D��D�|�"�[�(�ŀ$�I_��,v�G�V�{�K[/g�ȕSQ��TS\���9� w���&k���f�Ax	mV�O�BHp�o촁�[�c���C���~� �<>��d��$�paP�X�͉71C�v�������E��`���RC�PRd��Q�E��-���D��U<C��4�RPy8�����;o#�S��/9P�5��<h���x���[�w���%��������\��O��S��6��4�XZW��4��r���W�<�����Y:BÂuU�(W�zđ�+ް���Y���K1�{5]9��6�2ϠΆ`V�vQk���"ǔ��w��,�Juƅ�����mwj����K5xh�3��ǳT#j�x���DS�~��u�%�:�1�4�Ȫ��kR�����h�>��|y~}GDG�h(�7�=Qp�eS"��7�Nޱg��#͖��x�O���\p$�w�I����#u$����0z�3p������/®�3�ell�6T�®�b�f�6�!�-~i�ft>�B|v�Y�'�TE���w�2!���e3�B��V�<-��19�f�%'����՜�aGA�@�i��|�/��
��*���I��#�ͨ�=���6��&D��uU��r>�a����f̓������gZ�QE2�5#�D�=��oMO�	��+e����ǯ���S@3iT�^Ԡ���u����CX�[|��4�t���pzX��a��1�f`i��CZ� +<v�3�~��z��k�2���Y��NRs�e>7������R�q�P��ո/\��X�QG0Ƕ�K�葁�����.5��S���E��	ȩ��:D�r��J�~�U�����D[j̀Ep/cEwx]�Th'��Q{�-��A3�c�h�w8�!�6[���|���M�v��z�#����%",�E�K��׺ G��#�~�$��A(��@�Ptt�9;Y
���N��#*W!9�C�*ו���Oa|�����|�6<y�1 ��I���LO��7<z��g�4D�NB�O�~�o�Tt|�9�����x%8Ҩ~��I�����n�[�'=0�N#ڮ�ro2]���"�B�'��5.�HE��~�� P!���=d�}�D<������t����}��+�uu!e��:nט��o�-�n+�b'�ۥE�<����H�����s�J3��;�U�z��]@�0n��y��_�#~(�j	�0�sڮ�ɧ��nt���)Ƈ�M�3=Ծ1�eXI��u���\-u=S�꣹6� W/�e�QR��L�et�Uu��ψ��9?
 ~�Ym�?J�Q��^T �y�2���+�)��X��,��H5��Kl����W������i�������2��J��64>�0�T�@#$"!���>�|�����f_�E$�	Xx�fz�;z�caO��01z,�Qg)aH:�x�uX�>�I�z�3фbC�����&�F��fjL0U�n-������h��?��n�j{��L��F���ع�:G�W��l��i���|�m����n������&�a*�m@�S�a������~|�>^)G+d��~8M�9����=Q��)'h05R�$�:��TDl�>��b�Cœ����X��jW�L>�̕�Tj""����]{��u�Z�W@�ώZ��cF�Ur�J����9�K[���jAx�ث M���r��[Ԉj�XL���V�����&`�Sk���@q��aO�5�,�:(��K���:�9�,�gSd�K3q�����᫝Mgf��/� <�Þ|�/���2Dw1���wk�i����:����	&��:��/�T���+�f���	ڀ���☶�b�Ӂ"��l�Ж�&�
$��m�gi�)�$�Y)���Y��f����?�5 �k�2�Oڙ{��~M� <�-��R=���"��V��L����s�π2f
�Ҙ0�G�X���z�Ε�I��C�#\����W{���+m4��Md��İ�VmT��&c����j�;럞hث�L�W�Y&Z�tYw�iɂ�]�1Kh%��.�	6$��)�!Ǻ��EN�)7� _�q�G�?̤�,�E�r�4��C�)��Q-��2�xlnާ���w��:@��3����l9�]��܂��q�y��%E��7z�/Q�v��A>bW�.�`n�ޗd���1{�䌋(�8���֦�|%y��W� H���oa��h���b�Z���u�<;9.�������\$jDJ��7����������䅩��b�II�i��Ǥ>����T=�����e��l���	|!��7U�~)g
^�Yҕ_X94����M�pZ�䛍s��C���o+f5��M�B*]C�;�{ u_����4I��a�'� �p;�1��/��imI�{�x��3���?�:F����O�`	�IeQ 1�B��6�NR�u�أ����ח�a�?G��6��F�᧒P7�L��on�Wx�����OQ�#,���U��9�ں��� n��T��ܔߏv���`*���5�:�-���$/A�2��d��+}9�b�Xf�Q(:���0bȂ؅$��#KZ�>��s��Ң!T�8�LM��s��g���p�c�){����F g{�Р��\uh��:[��C9��� ��ޭ�$�7"�WH�w%'(a��ȋB�HE�Z�Q��K�1T��I嵸�i8�I!��5觢���W���\I��y�Ȅ���	e��k� xY� <�)�xWp+UIz��Ö��Cs��"�D\�xwJL�%X�0��}�@�Hdn�N�ء!V��v�`v0��*��g�B��Ħ��J�������cs<u�~E	�2�O���7���#]�L�����Gl��R�u���~Û`�2L��I���q>�U�A�j^?��q��юo᛻7��Lzi��Z�46)^�OZ&�V��z*7�p��Oԟ-�k fx=��E��1kؖ�6�BTy ѱV=_�t*8s�(��Hh݂���W���'~�-8�j,;����*m��T?ihc��;YnВ��<c9�z�t_$�~�G�y����Ū}K��]��Ր=ʑ���_���#�U ��TauXcS����T5"���{L�UG��܅f�:�����;�,:���zLe�A�u��g!�LS����0���©�R��m���1��}�}B2�'���9~!�?�U۪ܽ�c��+L%V�it�qf-M�D;��J �g� �\)��U�~o8g��\,=�Q��;�M�D�0_Gq�x��s0�h�/�1�W����Y�u�%�&�M��y~J9&�WB1�tO>��$�!.�����^��:#=^�4������UD����b#��}�cGذ�.�pN=�b�[�!��N�#��S��4����@����g�s�V�d����� 9g��:3��Y�<��j��]lrZY�&W�jH������9���rR�����Z���k!\�Ƒȯ�l �� �mT�l��>t�����Nv0N��W���e�Z�y6���8>���pj���G�"+�8�������PF+�v5�P�n��/�� $�w��N>.[����\a��=���Υ�Hm>H�n�E_��<G���t�����\��n�,���!�0�$s���Y�/�u�,u�"��mԴ=Rl��X��T5�U�/��jb��1�wS���4k�� ��G�ٗ�B_��[�*QV���G���!��9����@�p�0�����U�#S��4���@����Uc���D:< ƀ��Y���W;n�z�c0��$��~��A�˖�(�G�I�5�u<,�E�'p���_���
�wAy|�0�/�^!��b�1gA��I�jo�~�P�	#Q�^�tiI�(�7x��,ێ�Q# ,����=���5�_�hڟ	�t鎉�H�Q�*�ᗸ	Z��J����L�������d[�0��٠�W�̄ڔ�\ �757R��(.9�[��\�2��Q7b��?<D+VG���<��ZZ�3|��-�:r��"��	��ُw�&b��v��J>o�"h��o�FWs�����z��'�i�p��!����׺7Vq���dŸ�F�vX��=�������D���d�����b������	uJ�(Z�=�p���`�
��B#{4�9s�\%�]<�7�V���X ��zǣ�
f���Kq
�[������0"}1r#\%#����"i�.�\�ހ�n�p C�<��ᒤ1g�Js�t��H=d�-���:_���ܿ��3彆�{����L˟�N�<>��:�ĝ�Wq��&�>�ꚞ�q�ғE��q�jfĐ�y���ۙ�yC�΀��&ݖ�Ux����3����!��r[���x�D{��ͧ��+�����g�F߹�9��������A�V��&�c��i�ޤ�4M���\I�=%��V[��R�)��.?$��N�_w0���T�AC��j�an��#.C�V\�oi�糒�#��W�۪��cǍ�Z��pV�	h�m����T�ꮞhWk����-�������������a��zR��g��K_7�I�uJ�?;�$2.�uj���S
����)�g 
iw�|� S��X��?ѲN�>s��JJ6��&�6��Ь�|��"��(nۈ��^{#�u�^�e��0gn��; �{�Q>��o���d|�\}��q��8��^�-mqb^�@;��02{S$�,�f4�� ��Tɒ�W��rd��M:R�_'�s������ҳ%�>r�����5�!
\����s[�U���k��a���cH���$�R�^��X��3�51��a6%gvZy�� S�*+r4�|���V�Y`�o�ry�.���
������a����N~����6����F��LH�gǿ_����]4_Q.@��w�����.��p��oq<�@#�A�����h8EO36��~7���צ�h<N�M_ė�����f,/���7�[��z�}��
6�7�(�W��{�3%>h��B�]�ё�Tx.2f�L����L\�i=�6�.=�����1. ����+�d{M듆�L~��P���-Ed+�g;���<�Q���q�_����/`��Uݮ�0���!+m�:��̇�X �'��1s�	����ŧ�sK�R��*;D�L6�J��U*�a�"8�����y�k+8kdq��=/a	�p����{�8�r.��a�`4<@�+o}��Xa�L��u�X�=�u�q����ʓ ��!>s]ۇ�lӖ���yƏ�B`�}ދ��9�����}昶�Y���M۰8���Y�m����OE��C��0����%ԩϙ����Q���UX+��Z�:g��YoO!�,����������S�+4d�5�����*���;B#����xDo�hU��sQ�^!�7�[��b^�S+�M�O����s{����Kw�if;�D��(|�f��u��C��-�ݓ���=wٷ,��o�0��n���6��G�yc��y/�Sz�󛇆�ױoB��9t`�q���*ǡ���J#%*9���� �Vׇ��F<T+�B*����,	�E~���X|r�1���v�J�7ѥ⇩��LO�\��'@���[�"�:��p� �L�)g��/62����=j���=JBuŬ���7If��G�d�]ec��R@z�~�����yK�Fu��2p�־Hy���\_�>��8ڵňN?6��ԋ��ྂQ"�_d�E �ŹjdeI�3+Hw^�KK{�<�79�����Y��s��C�
-ex��17G,b{����b�RHj���_.���$e�c�BX]	E�����g��ZB밨���F�s)�מ�B(���'6��e,���A�9U�O~�nQ�?˜��QL0U�V��Q�ă2'o�a�QD/�\[�_�"i�"uyI ���m�a�&~�<��F���0�S�s�S�:iR���ΪJ�{Ӳ�{��Xև��zRZp8r�/�@d�ь�]U �����}�B4%Z��GgtGڌ�W$�KyrA�J�7��@c3��oy�گ�k��vJ�6\�]�_1���4�N:A9��_	]	���I�/7@�ؼ ��6�����?��(�o���@��w�C��֍Hd���zPo���S���0�e�c\h�BvDoؔ�w)�3�.�*���"	dH�w\�L��s{�3������Câ�^n#�W�C���T��?�|��'3��������U�!�0ʹیQ#DTr���dKw�R||H�KS��9�eu6f���G�� �`��R��bL�:������x@D*fK,�/���ʝU;��4�"���\��b�G�j�t�qƲD"̒�՜���Ù';��g7���Xx�ރ"|�,��k����}�ա_�|��A5���s��?H"��3�/��!�΁>�a�ʥK��X5f��q��Q*���7�FD�z� �L̫@��q��/6���H��8����M�����k]
�]�.{�o�B��5�f"`� &��:oLE���F��kϒ�fhh�������dt��f�-�$my���up���1B��
-��H6sX���<nً2>ni�S�z٫Q�Iϝ"������$�+vl���򫙎�Ru�`��cχ�	O�i+�G�hVn������B��<�{���Ӛ��	�����N���}16JR�n<ErUc-��z����0X��v�zs�N�1����Q�}��o�A�z�n�e���	����ƴ�5�Ѫ�{��8IG��u����<�T_y:�����O娺6��d!^xqIl�m�`��E��ݞd\�)m���
Q��H���S���{�%#�,4���I�����/2P^�/��U5�G�K��Gy-e�[�J�����ݪ`������8�
م�
96,�X��RG�Sd�7w5�N��4(�G�� ��:%۵b=*pOW�!w ٹ�ޣ�"]d�����Q�c�ޗ�Z�.�]t�!FH�ǣ�����/ �Z�ȸM�����E�����)H�(P׆$K���j��=�����=3SG�P6ŲPK,f�|�w�@3Os���tM��F\)��hئJ��:�h�AUqA�[;?��w!��Y>E;c��1�.���f01 (�N����P�[��CR��>�&1��������0>J�/<�)�����#C�D�.�������Ps�P��tq��&��.�"�c%v�I��+��ӄ��fd�p�Lw������5���~�w�Ut�\G9č���	r����T��f-�x$7����+k%.�0��z7�eJ���G�g��3�����W�b��JG_�h��+f�2F~�Mx1����,k�4�����F���>���;5~#%�~�2����`��zY$Fޯ�d��w����$#� u��o�������ƛ�T�NCM�M?<3���r����Jdk ~�f�YU���g��X��#͚���v����%O����6u�<�޾���_"nag��C�L�D��p!qL����Y؊J���	A�=�6t���`6FM�����L�z���ܵ�/�r�]o��p���g�:���\���f�oZl�M�6�C1�<9�x�y�T��K�g����K����Q���JU6�c6Ԡ2���s�ܖg!������E��*��Y�D�����drr�=iy����ڽ�ʚW,��@�-}��+���G1H-8M��V��s�J���R˅�m�(pQ#S4QD�;y�+�zQI��C/�l�P�	�LxO��x�v;7Ɣ~����j�������A�~5{�X}l@ݺ'�@� ���xf��aw�3w�j^`�4���M�]�%`�*2݁�憂���R�����0��$��?� lD�S�n"�����)o���6�B:���͋p�N��f�[�[i��s���1�B�^#�2v��e;V�,%x��y>0�ԁL\��E������U?!��
G��G��f;���j�����G+�h8[vL�pڟ�n�leBzzc�q�F"@	ʯ�㯼���4�s�Yo�AI�������E�~ey~PGL���R���^2���/ǦMٺ&��|ő��2YE;�㖅[�g�%�.�+?&��W2C]�����H��i]نNB�V������K��#
�ѡ��X�d$\�r����q�X���>0pV1{HIjpI�-�� �h��ƕ����#��g�r6�%�B)ѓh�`֟���h���ʾ]�'�Ɨ��t忥��J�*H���l^��:��@��Qn�u�۽J��5��@��a8��Ҁ̕��E�_WY� Ib2h��;�RJ���/.K�wA��ׅ��\(�סn����o�+��O;�36m�m<��&����0*�Ł]��S`wza�1����b�"���eG�Q�^�l��aG}~�=��a�^�� ;U]-K�����������v�9M%��<q\�fXR��[�D���GlC诸���ձs�1ɑ~,�ή����I��\���C�/D�3d�/8������"�������T@囉KG�(�VZ�������]Q�p�m5����
�ہ�_�G��� �d��U� �޸?����(K5����V����>T�\"�V�v���WI��PQ���֕��V�^��}�^i����'�����n�G]�K[4%"~�N p&{z��B�A�yM�]�~�i#�xR�C��,�<;PM�
@F�c����������]�S���\�U6������S��K�xF}���]���=�t�3�ߞ]���T(i�ե�?��h\~I���pım0ْ��Rfl
An�h������+��J	.��Y:UX�3.B��Љs�G"�G����q��lU>���\�|n	� ���6��}}m��v|����Q��-�s'/|��d;���TT�-�mG<~p2��ɥ����k���sǱԘ�2�����U��|uq�Fn�\�)=DҶ/�m�R(Es��=�ʣMN�K3]��"�
A����h&f�ٚ6�� �d��(MY��l9��*T�Sf��}��"�hl��1>��0���9$�G�(����¾b�=m�ZZ9���Qև��ʵAdK!�w�aGwD�Z-[��s�uӔ�c;��OL��qc�P�&�h�A�L䌋_4q���q�UR��3$keY�`�����_�ӻ�͓x7C����2�͵|D�Ŋrx�@zO���"[���i��Ms��zÂ���γ��1T�Z�]�qX7�j�HadS���]�cUm���<)#0�#Hr�<x@�*��W�@u����3���Y������ �;M��^9���!���T��c��(���t���m�=�I���Ng,O33$?[�����|l\�0�`=�!�N�_����슒���`��7ӊ��0�d��`e��B�]�O��\���@�cVj(���G���D�b�vrH��O�#�4���Iֿ�7 ��ݤ�����
c����Y@ٷa�h��1Z���FH�߽O�_TtX����!n�^�����.���N�QVq_9�ڻ����R��ػ���坋L�*������An�����,��q�4	�g�hY*����{9����6��C����x�L���f���ĵeY�wJ)��R�)�UQ�9S��@������^M*V@�	tp�E�JIR�8��G%I�g��C�l�͠�#��8�&X%3�s&���6:4.�ӑ�.���m�J��.,�!���&�N5�K"�Ē��8���"�������V+�]0�9�������^�HU��
��x%Ά�$[@S�~@�����o=��3%)s���W-E��PZ!��+���6t5�����Riо�]�t
�L�x�0�\��Cw2�qogl�Pk��ZAMwVC��J��`��Y���O�f$�i�p|��zvvI�mI	�Ou{�1�/Jr�ØrZݦӮ��nM �/��͙ҕ"䳵��x�CZ�c����k�J�@���|�P&֓��K6]~��%ˍ��P2I:���e����]�6�+�È�A�N:��+�yj1�c��!�LL4��`��t���1��i�fۆ�赀os�؝���
3*��� � 5�OG�k��M��Ny�(6���@=��1O)��2p�7�{*S�!��(˱��%��+�_W]p�?�E��5�\�5��w���'H�/Z`�Nr?3�ߕ�Y*0[��m�O�L��]7.�T��~��6�=Z��FP��TE�l�c5�r���X%u5%�.T�5Ǣ�_Hr-���������v����|C�w�Y�b�}Hs<L�-�A��TD�)>�Y���T��{5�x5� ��J�ۚ�C�p�ԩn4Dt�8U=�l��~}:@s��!0x���e��Qf�<�Z 0� �Ú���²Y���S}�����ibo!���OI��"F
n��l�>��9�mV�o/��&��G�J5^�lpClngsS8�W���H�Q<��D!�z=���/ Rj�Vl�����䣤�)7�����Ǎ>N6#��ߜ)��Y�(W�lA&�`���NZzѫ+��}~'�Y[��<��O�:s��V�Za]	q:]id/����:i>Y�L�h�Ү��m@��o�U�=6%h=fyۀ�xر���zQ�H���x���|��mH;������P���{��-�1~2x͵�(���6M���-R ��"]W��5ު�i�$��ףb�w3�|�N���m�y���h���퍉���p/N����_g㾯;Y�d]~Q�&��WKrHO��\+��
�֜���e2k�,�#���@g��$��q�w<��2CB�HM�&��M�GaC@B�[��y�2ޝ�(X�<������e��΋�w���]��F�s����N�9�6�ZF��?b�-��]|�l�N��Vσ�y���Re��4���G }�r� ���U
�6�3gV��wKH�}�^�s)3]�g�/(���g�.�1�}<؀�9� �����̌�h�T;Z����>��gwf���E)�t���7��������8%���旍���4g��XƆ��'eK��B����[�m�nmP�O	0B�_����uҍWhg����f�|�,H�Cz8 戱�����b'������̶� ��˃�kҴ��V������+Xɸ	����LX�����5a�W�?�����z>�&�xO^d�i�����8���ǵ�����PW�Rz��c�%`���kh�Q�a�S��6Kq��@Z�&b�в$I�ߕ�S?�'�z�⊞�� ��뱶S.+"̢�|O�|)Zu�. q+�4?Y*��'i}6��7�/�R���S�fN�P3qS�-]*m�J�O��|��Ɲ�Z�T���L[Xf����zMs�;�\����7r�-�@�>zly� ����4m�Xn�?���F��D��l�p���K&�h 0��;J/����q�	/��0,�/����h��>1=�2�����J�cy���}�w������H0*.5]V��B��Ɲ5,���>ר�y�Hꕽ­�)�o����Ί@�^A�Ӽ<��3��rZ�h:u?ŗ���� ���J�?�0T��_.���Ǣ�TP�U(P��*�߇JP�m�&g��e��vF�9^%C���#xz���'U���
��vo�f>�0��	L n2�J�;,�p�F�^����rzӰH��6
R�C��V��m'¢�2��%���o��&JP`5��X�l�:��<w/̄�x]�#;�񄘤5BF�%H�ن�IW����H����R��Ta.�lR��MŃ�x�&tے���mB���qS���kt����J2\����3�0��
=?9`}8~�㽙�y�~
lZ�&���\��W��;Z%�,����z���5*�LV5صj{��֒R�����[�Z�K��鰖��>1��v�WMGHI���\]8J���V�b�	��|�n(ñZ�x���A.d�̗��r*d��Ol����Z�zO@y��
��2���X��Q����]]kE����T-���xƲNþ���b�T�g�����a�@��g�N�_�8��Z�F�e�i�%����e>�0H9�B�R��+u8B�6��Z�Ym���Wb�a>�"Mn�0�d��'QF�_��ܚ��"ڱ4�幰�;��凹w�2m�S�y�K�f<�y�vs*�V�WF�'(F����ua���`p���
�~K�l��Ig	��%vn�Ub��`���5S���T��`ג68)Y���KG�7f���T�d�ۆ��915�oB���hR���y\�HVoŨmLJ�vc��$�3G��!��A+���0�^�=,	�Vb͕�3����NG=��U	@�~��������d��3�ಏK܊��X]�B6����k{_gE�T^���,�"F�m�d�q�e,�}+�|�U�x��8Ef��,.�3q���gt�*Tg4ߘ�1@����;d�+��
	���~�E(L�/�G�r.�т����}`�� �8��I~�Y�_�kT�B�͖������IM]�@��ҹb�"�ޣ�e�b��\��R����ы:����'n�ҘK��Z�>�{D�w����<;a�^ O�O�P�G��1�=>�h���	��t�&L�8\��\�����L RZZ�K~�u3Y�/�粪�Od�^�J n �ڨ�{�n_a�J������o�Nw��*� �,X�+<_��~<����%��41�'�A������kh��8�Z��vg��8�B3iS� ��Ex�iq�vA&�^�E��DW�ЙH�L��\��^V��|CǞ�O3�q�-�Bu�>R�^��\�_�rjD�;ݜ{T$)\>�Vapd�{���O��'�G��e�����k
�e#�*r(ѿX�閧��i
I�SeE3Cfi_n7������-����.�s��'�l+4wȚ׾��M7��*�B�q�7&���}XaX"����Y���:Eh�����:|_������&��o0߬vj|���Ќ�!��h�bÁ�l�kW	��zXÊ�ys�_� �]�]���C��khd�X[�O�)'����Fa8�����t�0ޯ��kY.�m'8ZR�sP�/�N�3:���h@/}2��?�,.�^6J�� �Y(��s�6��}'D��A������J6�P�g_Ј���X�*��_�y�=ȑ^�<�&�� �?P$)�xN2'�K(�8q��x�����\2���i�9{�A.E�x����kP��qï��sQ�X|�q��<����sA;b�Łu°�1���Z�q���CO��X�U�K�f�w&v%�s t�x�kl�WF].c���ۧ�K9�8�� ��T� P���CI�{�36F!�9V	z8�5�R�T6��$ݩ�5��[۷�)l�'����kȁ^��V�(�+��m��$T�՚�Q�'��G�xC���ގyl���l���[���rۘ��k�eXh�+o2�[�([]���������:����=e�p�y�%髦�Z�4�
�ޢ�O쩝�� L ��� ���e@�%�O?F-98~�@�se5k��Y����n.lUx:����@��3���t�=$JP�ƄV	6��T'��x���iQ�v:]��>���nB#x�J|ҳg��e!8b[��鳥�fHL�Ew�ɺ��W�=��QU��H(S�f�A�~sã��kWz�c����M�L"��*�όs��.V�W�]?`KL�x��]�yMjrPr�c���L
V'nz���������)S�%�t^�t5^a������b��0��� ,�Y�v4O��DCS��S����w�\F3k)d�}u�~ʻ_e�^�+IH�׬���a�@kS�
�K������L������<�P��U��ɁP��0��u�K���C�%��ڂ�DA55X�׬ aX$��c3x��3�j�06�4��{>}Q|�����H��d]وn�V���h�f����T��:�>̭�X�eNWn��0 ��l�������0 �Q���Q!��h�©rݬ,��0�˵�H�J"�T{�~��v渨�ތ:�<jY~AW[e�Ր98�K �T0�
O}wW@J����z����16|��fV�=�ϵ�X��E���0K�FIe@B����>�i���5x!�OhVU�n��5^����{�xv�$��DurYV�t|�!E��+�qK�r���Ϯhu�`7!J?��B����z*4�D�iG�k�g�ȵ[�U�^�G����F4qћ8���T�6�΋0�52 w��|�� �Ѓ4�������b�s�|�'l��Y�MP�~0�^����H1�g2���E�dEM�vmꐖ$�R�=/��+fw>���]����H`EU��9 �a�5��)J���y���H	�gw�W1�2�ݧ����O��
V�����p9�'I�FU�r�V0'%-��xv���;怜��-���;5��J�����RBNLhqE_VhdYu���B���V�*Q���C�Ӝ/E�]A'�P۲	1zK��h	QR�H��W���6�fuä�E�6����Ce,ƺKRlaQ��h�
51N���x�,�4�=���b�>��k������Ǣ�T�HH�v�����gfNٝ�������^����i�J��g��!"%�a�6��_�\�Ś�%�M�S?`�`���N]T�Kj��8�U	+�eO~Y�V���أ�/A��ra�Y�Le�`(6|aO�����H�V%���h5f7@�<n�>� �f��,�a��#���x���:�$���AZw~y�2o�T��r�c�c��e��o�m��
�P��p��}��cO�I�»VV�����
#&��J��P%Ne�4�Ô���b\ήܣ��ɹ}YH�\c��xC�l|ʳ���KVU��cM�=O�={�1��RT*a��N$��^{K	�������4ґ��q$�ع�Jܝ� �j�>���>d��xHOQuIm�tca�E�ÆTJ�ɵ�`�q��s���ؼ��S+��<��J���1J��ToL�9�j�j�>�<u�3q���F���Oy�k΍�7��zPy��#����>^��,R0��飄F�bH.5���O�@���/(�
-x��d���$�T�ژs�����k׳ܵ��˃��\�<F1��#¾���?H,H_g����zB_��K�Z�0����Eߌ��i �n����P�q���d���,����z$_҇�)!W�T��oMc��E`� �Y����=���OT^����./��󲓒��4Z�)&6���7�ޱ������.y^��:[�>��3�Wa�|MڍN�+_{G\1�'��D<γ�<[��4]� �p(V��c}�� eN��ē]�y��(g�\!q0NQɃZ�����V',��X���FwP��[5d+mѯ#�mS �R%y��4Kѯ%\g��NT;M,d#���Y&ȵ�q���t���$Zew�5c�ܩ��JLQ���G5���]�:��",mԞR��ِ��.rJ�D�f�u X�s"`7{���ث��yK3-VM�,�OǊ!��4Q��*�A�7���~z�nz�������7�D��y�8>ԯ��>wv��<X��7�@�+�����FכBAmqD8&իΦ<#f��m"��-kL�T㶗�-�@��e>�Zmey����ͷ�
�����[�l{��r��)���e�d�uG���E�I��Q��Q0�>J��t�`��:��]OM�4W��3����-�=5uW�%��Kʌp7�?�ꨋp��;2�E�v��Jf�2j��84��ЕU�Q�k�[�<ך$���h�_<T�D�9��'J�`fd��'���L#{P
�H��׳/4�''d�{��$���^�|�E�C+���R�ϞE6���
1:#���T.V�%�Tķ� ���"UW�klӕQ9L�?�� {���)��}%p`;0h#|fӰ; �yٟo�.Z��B8�S���p�1�����K��x ٘�+��y�j����t� ��\1h�����^i"#����|d�i5,q����?�v"�z�G��C	�~�=���
��s�h�4Eu:����;E�us����?ZL����K�5Ɠ�E}�_9����A�ѹh���c?B�'I>TzR�uù��_��g�2�
��-�`b�gl�i��%�{𪶅��",��P:�fX`�[5\W6����j9�!ID�c�[UR>[�5�M�.��}�
����\��Ǣ���1���9�xLQ+�'Fѳ���|��"�6���ի���AR�'�?SR�:��3~�V�ul��+E>�x�
�{�J ԇ ���h6�fнpm,�G��)�FZ:2C��|�9o"��A8�џ�JJ���t�� �Mr���#�a%�p�t�r�w}�WҎ���bA�g�Ş�*;n�`}�E���a��`�L����Pụ�nE�sa�\��y:I����qsD�x��V,����d
�FP��p��rw݇���w�}j0�����F����Fa�nI=�x�ort~����@�cn��|�اcǾ���s7�o���^�m�$i\̺E�J�l^"��*U�A��%��[�y��pD���]7�[�܄qmƞ(��S�\u�l)���Qu^Qϖ,;z6�,��ж�Ń��?�V�<?|��Sv��9�����%S��zB����@�&ں��-q)��Fֳ������D2+YR��A��n�:O��RX䳶'� @��¢�s��8�d_�խ���(<I�b!�T�6��p��=I$�#eb$M�ALp�m裣B4Eѡi�b�8��:�/4���w��}��-7_�'���A(Ц��[@2�EX2��%�� �aU�n+�k��S?Ó
���m�����Q�]Sn��?���OY_�+�(�.��	�W��~��\@jf�X�X�˛3�mT��%$~�Bռ�2�b��x�$�B����4�� GËӠ��v���������*E��@|�J��=�;�ϟμ���5d��d��q,j�q���ߊ���,(=�܄�fY�2�n��8��,<[�p5�z�wQ/ئ�ұƋ{�q�oz�&O�W{d��+�j��>�9�\�<�lz!�Ĝ>M�=����/h�xp��)!gEg�[���i��ş�v�C1C'���"�S�26d@��MY��ʔ�L\���r��}^A�F��q��-�WW|�MB��������Z��7dڊ=��������x�UiNu�)D-Y����ͤ�yԮ QB�"��B���NZ����)�U��� ��)���,��i{nڟ�822�8Մq�p���`Za�5�"ង��.m����n�塋!����ƀ(��"��u��ļ�����N���R�|<�E8��}��e���Y�c��AGe��2�x߭���YҩH���j�+o�{Z�QB�HkINV���P���w%�?z�ݳ9��`�5�����2j�~e0[> ���p.�;3�q�/��A��k�.�ZĶ)���~��L��q��]܆Ӡ���F��o�.蒜���`�s����½��� �q{���Ǣ�cnM]=�3쓛��<c�[���}�p�|��%�u��=�p��CЖK�Ϭ�%������]½�C�o�X�^�iDq�Hr	��G�E<1k'�N`)�`��+�%ѝ���� _�ʧ5�w�wn,��Y\R�D�4���&�(.x�������CC0#g��lAxf���c�T>�&���C_�����i��j�=�[�y/��
��_*���u��'`N֩f��ta���������WA-����m�p��T|�z�^s�K����U��|��	�ZLD��~`mt�R��+���F��!��ӱoͻnyÀ�L��HV���8��2�*D�u. J����N�׌��Τ����}P&�W�@8vp�:�7<<@�֧�+�hopi�v�p�K�!Gnn�uhdA�?�°�!�ҰY}n���a8�GF��9i]�Z�5�f�P��l���"ˠ����&�@�6;�F�5'���P�3�W��kl;�����t@�.E��wy�{��*��ny��*�9�qb�b�<�{c� doǲ��H�����n���6|�T�vU�b ����q��y4{�(�lU��vCK'�?Z����q;x�~��s���=��F�ay{������"2+��3�^�S�������/_?��p��Pu�;�D�d�ԖR�1�4Í��K���6i����:\�e��>4��*)4��y[JjK�Fz%;v:u<
��eM���T8u�M�����=�Րo�4Ґ:o#�+*�6��k�M����"MiI�K�����3��}Y��[��F��s���}<�W`|?�Vb!�C��n�u
�~���"�Ң�
}Pճ���ʘ�Zi�)M���Y���aG#k9A���^��B���|��u�A�0�m��x��IDչ�.�����Y�NvY�����?�N�U��l\�K���vWh�J�T��^��usW�%+��?S̅o�]�¤Ǝ�c�9 |eZ�r��GƋ��J�,����ނ����CZ����rqKi퇚��a��Q��?��^��_ڑZ��Ό���J_;_�!�Y�Iqa���1�P�K�IX�\Ý6�������3��_k�#�q��	���q���z0{�T��q8J�����T�C�1J�$v7���򤧝�B��QQtW{+�mە��Pa;����sJptn�"�a�Ph����l�˔�|~QD�\,0��mHEs������`V�1M�ڞn6��<�C�ͥ���ie��S�ph:�l�<�38?%��{�z!�~e?+�L�6�^�\p�߹�i�����0�DJG��%�B�ek�g�<�:������FT��y�tC�2���6S��iK�~��z)��#���NL�|^�9�sT�����Y7:���N�ägB�dQ���g�]B����������v��ږxJa[�c�����gIU��x��R����jz��|���5��Q�rXVһ�Ed'��h��#j�ƹ�ҫ;�X�IN���Rq��ܖ�z5w��ٽgF�rz�"Fs�U��~0��"mf�܆ES;%M��|$�$���N�:*']l*Y�Ij��B�7�TmDP"�E���co��Xߌ�W�~\._$�{;������UN�������Vl1�U�
'�%m����ݨ�@�*�y�f!�O*
G��S'n�}�ܦ�h�a�	�&Ë�)���]82��fZ�7��c�0q]�G<�O�L-I�K�y/�P&X�p�}'��,)��+c��t	pz}s���Q�U�g�Q0��WeTSlUT|�eo�.׶��֮��7'���W��?L#�&��z���ۻ����Z����%��G"u-m���<�Po"�K��]J���v�K-�P&���;��R��N�
ݜ;<�g���"S5�/:�A�r�W��G�oyl���@2���(�-)S��YF�L.�ꂙ��T
/p�1 /-��~�L�����	!�Il�:/�j���à�t��Ƅ'bP/]���`H�Ow|��%d���e.V�Y���=�@w�jo�Jdl-�w�,�E�M�5ɚ����%M��Zt*);�!E��w��
uȿ�tj�$�IHQju; 'Ơ5���ٝ�^i�:�n�Α]h;�t��t���;���&C�ک��4�ܕ����8f�.�!)[�%�{�u��m�hD��%�o�ZPB=�]��m4�ד�������̳��U5��^�vFI��֦����dU��z؂+���Q.^�*�3��|\f����I�}�a��R�PEٓ����1��M�5���/l1$�������J�
�Gq�w�oS��]p+0ph��� a�����������0����z��ɒ��G3�Pɩ�D�@��aa���CW�Q���C*	%���� :����
zՠ]�6*c:'�n�C��|�Ly���-���</T���7�\Q�b��G$q\:�ww�� \�̇RIkQw��Z��L?&�����M���z��,����Q�E�@F6�a�j���J>���o��o?�i�UȒ�����v*�~�*�a(0�;��f�٠����[Fc!L��=��o���exiiR��K�v�K?�ЩV8�3Fn��].,��RLҗ���A�ߒ۟E��#R��pY�g��렗hS<����t�W��MI�)�����%ͻ�Bs*���<|���L��vU6�{�@�MZ�a�K;���u}WP�C�����h����J$	D?�?�@(��t*���Q�Po��l��P�=ج�ϒ�N��,B=V�x��0{��~��=ڷf�	�oJӧ���U�@�Z��ͤ֓���[T0���QLr��l`!���� ]UV�.���2���1C�6�{��)&Wܳ7�����B����4������D;��Dܵ�h4��j�w#N<�!4Z-���ؑ#�p�ʍ��s�[S��C��j��L����vK0t�,�/kG;L�?(��=6H<�j�ƫ޷��L@��f��N�im;�x�H�BjzC;ゆ�g_�=`�ڄY�*�����Rv�]��$S��j/�'Ue�(B_�������gm����^����rz��n�8���7'&�k D�)�)�BB�b8A��Y�uD��"$F-�r�]5����FAd�?#݂�!�nP���6F5��R��A}7&���Q�">A��@���Ԣ<�E��}�媒e]���9K|��3��k�{��z1 >x<�J�
��Q�Vfk����ў�1��S�v�4'���ڀ�MR����c�����Z,uzļ}�^M=������ ��+���KPnU��7�{�1�o~.ӗW��Ċ;�dUX����D�$-M����S2�2u���̽��1�S)�
�ۭ֘��̂�����V�*�q��=�KU6;p�������D,~��>7��|�1<)�<+�W�	V�H��P���c���hd��f�qc�Y�\�;��1���j	;��|�_p'[�lF$g�sM��S?$��L��.�?���o��hK�s�8��Wq���Sv�O��(����|�6�W�#�p3����0���&2k���� Y�+��I��R�����2A`H�ԑMW(TB�j^�{��Wh���!�yQ�G	,�%�z�懠J×����m�s4p"j��y�X���Z\��vMTI���/�^�מ����m{��Ӳ����P.��v��;=H���΀�|�o"����=���� d����bk���ɇ��⃌�����&$�(�?<���f�{y	|����SG�IgQ�&%��t�2�g���D�&s��Z،�X_
�����r�In5 y<�٦AMJ�o���/��K�]I�T�5�uW����,�E�+��0��uǇ񧹼�ޤ�D�$C�L�X
4C�i��C���=f�j'o��r���.�ɁAփ����h���� J�(�|�Lx^l�ߊ&R��i&���7+Z�7�����]�v�,��{a���"z,qr�mh�2�S��n�O�` ����'(C- �Zl��Xy.H3ڧ���.��`�H�o=[I�ua4���K�N/ZvǬ�#X-����wi�ۂ��F��Pk`>�ž`�#�pL�;`�X#�7���v 9�Ē"�I��y�ұ����«OH������Mc���K[^H
^5%�omPV%^�"�esz��/�M<�'ՙ�Ӑ�mj=o*̘a�ax��[h��*���'ZR�/&Xx�&w�/��e�;.Z=c�$�2����(�m�����
�� ڭa��������W�{E-��@�n,m��Z�"h�������V�-�J�K8�F�O�"���L)�>�t7K���Br��@I\%�yo#h�
X�]p��;F.3�XUG�ڎ.t9��'�t�i�jV�(���dh�p��mK"�EʹQ����P���m��,�zX��>��e\ˍy�)L���l�̉rH^]%�U���2K�B*��:R��ɭ	�1��RBbuX�u��h�
U˶�M�P��ڪo�Svw��fS�H���qኅ��B)�����=v́�]�3�6fj�~��l�e�"��=��9e��Xʃ��>�De����i8���$�V#;O��U���0��죅s>."ج7"G��֋�������U��F,�/f�A6w�p���F-5\,�	�sR~�kvZ��kI��ޤ�����dM������X�ي�� Qi�pDvӣ^=�=J�`{�:H@eJ��s�	�i�S��W�y`p���� �/뽬9�W<�]:��M=���S�V��l����T�_Ց�:_��UH BC
�_�oJ���"|3��5s���%�e�TY��fc�V���0O�ո�T��.���m�������ҧŐ��>�!F��#^���&�x�	��R����xoW?!�7F-�5%�s���:�u͹7�{&J�_%e����(Z�!u7�����S��
V��gNB0�=I���q���$��͠��b�m�U��ɍ�P�� ���s�� ~X�d�I� �	y�V���_6'����憛��Ʀhc_릏*aiCȦz��G3��A��fgR8�BSG?���Zʧm�t4u��5��$7Ԗ���54���"=T�Iy�L�}F��HP�-����p�X�$���I`����G"<��$�U|���۸Io��*唗��w�d�W��@���-?D��|*M�g��Ȑ����(~�T.u�}�J��*�jȦ.�Sq�y@�V�[$D��fӔd�%�Uj��>���<�v�����@mm��!{P�T�O� ^�!��[)`,J�G�.��*|�L�M��Z�ў ovV�ƻ:q�\�"�y-_������#��8DR!uڣ"}M:f�;zD�0jI���P]ةK�h��MQ=���QGSD7���l���^L�.B^D�7�	���J�c	������a:�-�&�o�&~ȋ�%���1���Ce�L:2��>tPY3���_�\�XL)�3g����E�!���	ā{�13�<���D6�u�ߥ�.^߭$ӡּ\��J�%�Xe�QK������u6̓Q~߆V�aD�������5�V�F�i���`p����Ass��&��Y�]���=s�zP�bC���r��.�
=P��eYc"c~�����ڳ��MP� ?d�����gu|1@7B��`�!�>R_�CF��X�(g��$G�w�����#��6�Q�Dަ�y>��p��ȓ�-B>*bJȿ۹��/]/�q�
NӲ����B�&�N��Sw�����7�9�6n,jZ����$�D�gP7/�7Ab�:���M�xS�[��j���	��ڍ̣����Y�`��� S\ll�l8���-:ow� �[����������"��͞��9����O�s֕{�oU�	�e�� ��%?(�y�c�\.�̚VQ�!"ޒO:��R�D���DO�M�)��*y_8�2���F\ӲN�-+���su(ol�����ɾVD$�pj{Xۮ�q��h�v��Z���H� ��r�0�܍M��Z�W��+�R|�.�j����e�dϷ�%oB9*��\���xc�@�$��L�q)��9V����+Y���U�
�f����/��H��"���4Y� a�UZ������+�W�CN���i	ڧ,��
�2g��d��!E��ljB_R*���I4nʏ�ht����	\<������,�{�$����S���nQ?=�����;�awR!�W�V�n\���C&u�f�+|��LC���+���5��b�7g˝"����DO!�"	���Rf�D-�k�<t�n��j��.�&����;�,J�\x2VM�V~3�K�.����c�\�&�ʜ{r"��s��w��P����_��J���Ff�F%p|Hʬ�]��_n��q��ߥ e��iT����b��-�)��������9�[7����i/e���a��H�(��H����w�aɉ�!�wGN��K+�'���YJe��k���@�0��a[+�d��ϙȞdT�N#���Ϲ�x��=�����@Г���w���Cr���z�\@�$U(uz���~�@t�	K��Z_��Y�8��!��_�����6�)P�lgġ�&��[�	W%�K��Z&�:�;����ʉ=y����ω��q��X~����Ԓ��M�6�_��$��1��	���� �^�$��8���8�3����	Ŷ�|v���nj�ojb��hY���-��3�.@J��0')cܻ�sT�n��N7��sy�c�W}>}�M���~�bې��=�{���v��'wƵ���r�t�F�8\���t1��:��9t�Tv�|���Gm�N
J��bHk�